* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__nor3_1.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__nor3_1 A B C VDD Y VSS
X0 Y A VSS VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=17000,540 d=9350,280
X1 Y C VSS VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=9350,280 d=17000,540
X2 a_1390_720# A VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
**devattr s=34000,880 d=18700,450
X3 VSS B Y VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X4 Y C a_1560_720# VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=34000,880
X5 a_1560_720# B a_1390_720# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
C0 A VDD 0.11749f
C1 A Y 0.08442f
C2 a_1560_720# Y 0.02841f
C3 B A 0.06746f
C4 a_1390_720# Y 0.02048f
C5 C VDD 0.11645f
C6 C Y 0.31843f
C7 B C 0.19861f
C8 VDD Y 0.1637f
C9 B VDD 0.08472f
C10 B Y 0.14221f
C11 Y VSS 0.51473f
C12 C VSS 0.3391f
C13 B VSS 0.33074f
C14 A VSS 0.41565f
C15 VDD VSS 1.75446f
.ends

