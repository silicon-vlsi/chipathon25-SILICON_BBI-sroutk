** sch_path: /foss/designs/work/xschem/gf180mcu_osu_sc_gp9t3v3__and3_2.sch
**.subckt gf180mcu_osu_sc_gp9t3v3__and3_2 A B Y C
*.ipin A
*.ipin B
*.opin Y
*.ipin C
X1 net1 A VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X0 net1 B VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X2 net1 A net2 GND nfet_03v3 w=0.85u l=0.3u m=1
X3 net2 B net3 GND nfet_03v3 w=0.85u l=0.3u m=1
X4 Y net1 VDD VDD pfet_03v3 w=1.7u l=0.3u m=2
X5 Y net1 GND GND nfet_03v3 w=0.85u l=0.3u m=2
X6 net1 C VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X7 net3 C GND GND nfet_03v3 w=0.85u l=0.3u m=1
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
