** sch_path: /foss/designs/work/xschem/TBgf180mcu_osu_sc_gp12t3v3_and3_1.sch
**.subckt TBgf180mcu_osu_sc_gp12t3v3_and3_1
**** begin user architecture code



.INCLUDE gf180mcu_osu_sc_gp12t3v3_and3_1.spice

**Netlist
Xand A B Y C gf180mcu_osu_sc_gp12t3v3_and3_1
Cload	Y	GND	10f

**Source
Vdc	VDD	GND	3.3
VinA	A	GND	0 PULSE(0 3.3 0n 1p 1p 10n 20n)
VinB	B	GND	0 PULSE(0 3.3 2n 1p 1p 20n 40n)
VinC	C	GND	0 PULSE(0 3.3 4n 1p 1p 50n 100n)

** Rise/Fall 10-90%
.MEASURE TRAN tr1090 TRIG v(Y) VAL='0.1*3.3' RISE=1 TARG v(Y) VAL='0.9*3.3' RISE=1
.MEASURE TRAN tf9010 TRIG v(Y) VAL='0.9*3.3' FALL=1 TARG v(Y) VAL='0.1*3.3' FALL=1

** Delay Rise Fall
.MEASURE TRAN tdrise TRIG v(A)  VAL='0.5*3.3' RISE=1 TARG v(Y) VAL='0.5*3.3' RISE=1
.MEASURE TRAN tdfall TRIG v(A)  VAL='0.5*3.3' FALL=1 TARG v(Y) VAL='0.5*3.3' FALL=1

.MEASURE TRAN tdrise TRIG v(B)  VAL='0.5*3.3' RISE=1 TARG v(Y) VAL='0.5*3.3' RISE=1
.MEASURE TRAN tdfall TRIG v(B)  VAL='0.5*3.3' FALL=1 TARG v(Y) VAL='0.5*3.3' FALL=1

.MEASURE TRAN tdrise TRIG v(C)  VAL='0.5*3.3' RISE=1 TARG v(Y) VAL='0.5*3.3' RISE=1
.MEASURE TRAN tdfall TRIG v(C)  VAL='0.5*3.3' FALL=1 TARG v(Y) VAL='0.5*3.3' FALL=1

.control
save all
op
tran 0.5p 150n
.endc



.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends
.end
