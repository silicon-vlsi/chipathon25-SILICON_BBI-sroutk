** sch_path: /foss/designs/work/xschem/gf180mcu_osu_sc_gp12t3v3_and3_1.sch
.subckt gf180mcu_osu_sc_gp12t3v3_and3_1 A B Y C
*.PININFO A:I B:I Y:O C:I
X1 net1 A VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X0 net1 B VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X2 net1 A net2 GND nfet_03v3 w=0.85u l=0.3u m=1
X3 net2 B net3 GND nfet_03v3 w=0.85u l=0.3u m=1
X4 Y net1 VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X5 Y net1 GND GND nfet_03v3 w=0.85u l=0.3u m=1
X6 net3 C GND GND nfet_03v3 w=0.85u l=0.3u m=1
X7 net1 C VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
.ends
.GLOBAL VDD
.GLOBAL GND
