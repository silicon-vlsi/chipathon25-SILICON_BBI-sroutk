* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__and3_2.ext - technology: gf180mcuD

X0 Y net1 VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.561p ps=2.7u w=1.7u l=0.3u
X1 net1 B VDD VDD pfet_03v3 ad=0.62333p pd=3u as=0.561p ps=2.7u w=1.7u l=0.3u
X2 Y net1 VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.31167p ps=1.86667u w=0.85u l=0.3u
X3 net3 B net2 VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X4 VDD net1 Y VDD pfet_03v3 ad=0.561p pd=2.7u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5 VDD C net1 VDD pfet_03v3 ad=0.561p pd=2.7u as=0.62333p ps=3u w=1.7u l=0.3u
X6 VDD A net1 VDD pfet_03v3 ad=0.561p pd=2.7u as=0.62333p ps=3u w=1.7u l=0.3u
X7 VSS net1 Y VSS nfet_03v3 ad=0.31167p pd=1.86667u as=0.23375p ps=1.4u w=0.85u l=0.3u
X8 VSS C net3 VSS nfet_03v3 ad=0.31167p pd=1.86667u as=0.23375p ps=1.4u w=0.85u l=0.3u
X9 net2 A net1 VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.4675p ps=2.8u w=0.85u l=0.3u
C0 C VDD 0.08642f
C1 B net3 0.00871f
C2 Y net2 0
C3 C A 0
C4 net2 A 0.00375f
C5 net1 net3 0.00169f
C6 Y VDD 0.18192f
C7 Y A 0
C8 VDD A 0.12462f
C9 B C 0.09692f
C10 B net2 0.00375f
C11 C net1 0.14156f
C12 Y B 0.0024f
C13 net1 net2 0.08029f
C14 B VDD 0.11714f
C15 B A 0.06819f
C16 Y net1 0.28319f
C17 net1 VDD 0.6672f
C18 net1 A 0.22916f
C19 C net3 0.02615f
C20 net2 net3 0.05362f
C21 Y net3 0.0087f
C22 B net1 0.1824f
C23 Y C 0.03198f
C24 net3 VSS 0.08046f
C25 net2 VSS 0.04401f
C26 Y VSS 0.31276f
C27 net1 VSS 0.83934f
C28 C VSS 0.32317f
C29 B VSS 0.28589f
C30 A VSS 0.34197f
C31 VDD VSS 2.49623f
