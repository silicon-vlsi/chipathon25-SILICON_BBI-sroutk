VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp12t3v3__nand3_1
  CLASS CORE ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__nand3_1 ;
  ORIGIN 0.850 0.000 ;
  SIZE 3.900 BY 8.300 ;
  SYMMETRY XY ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT -0.100 4.550 0.300 4.950 ;
      LAYER Metal2 ;
        RECT -0.100 4.550 0.300 4.950 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 2.800 1.000 2.850 ;
        RECT 0.600 2.500 1.200 2.800 ;
        RECT 0.600 2.450 1.000 2.500 ;
      LAYER Metal2 ;
        RECT 0.600 2.450 1.000 2.850 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 2.210000 ;
    PORT
      LAYER Metal1 ;
        RECT -0.300 5.450 -0.050 7.250 ;
        RECT 1.400 5.450 1.650 7.250 ;
        RECT -0.300 5.200 1.750 5.450 ;
        RECT 1.250 5.000 1.750 5.200 ;
        RECT 1.400 3.500 1.650 5.000 ;
        RECT -0.300 3.250 1.650 3.500 ;
        RECT -0.300 1.050 -0.050 3.250 ;
      LAYER Metal2 ;
        RECT 1.300 5.050 1.700 5.450 ;
    END
  END Y
  PIN C
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.000 3.650 2.400 4.050 ;
      LAYER Metal2 ;
        RECT 2.000 3.650 2.400 4.050 ;
    END
  END C
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.850 4.150 3.050 8.300 ;
      LAYER Metal1 ;
        RECT -0.850 7.600 3.050 8.300 ;
        RECT 0.550 6.250 0.800 7.600 ;
        RECT 2.250 5.550 2.500 7.600 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT -0.850 0.000 3.050 0.700 ;
    END
  END VSS
END gf180mcu_osu_sc_gp12t3v3__nand3_1
END LIBRARY

