* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__nand3_1.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp12t3v3__nand3_1 A B Y C VDD VSS
X0 VDD A Y VDD pfet_03v3 ad=0.595p pd=2.96667u as=0.595p ps=2.96667u w=1.7u l=0.3u
**devattr s=34000,880 d=18700,450
X1 Y B VDD VDD pfet_03v3 ad=0.595p pd=2.96667u as=0.595p ps=2.96667u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X2 a_250_210# B a_80_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X3 VDD C Y VDD pfet_03v3 ad=0.595p pd=2.96667u as=0.595p ps=2.96667u w=1.7u l=0.3u
**devattr s=18700,450 d=34000,880
X4 VSS C a_250_210# VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=17000,540
X5 a_80_210# A Y VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
**devattr s=17000,540 d=9350,280
C0 Y C 0.12513f
C1 A B 0.1103f
C2 VDD C 0.21445f
C3 VDD Y 0.49739f
C4 B C 0.09637f
C5 Y B 0.13088f
C6 VDD B 0.17995f
C7 Y A 0.2013f
C8 VDD A 0.23323f
C9 Y VSS 0.50813f
C10 C VSS 0.5083f
C11 B VSS 0.4242f
C12 A VSS 0.45023f
C13 VDD VSS 2.23521f
.ends

