** sch_path: /foss/designs/work/xschem/gf180mcu_osu_sc_gp12t3v3__nor3_1.sch
.subckt gf180mcu_osu_sc_gp12t3v3__nor3_1 A B Y C
*.PININFO A:I B:I Y:O C:I
X1 net1 A VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X0 net2 B net1 VDD pfet_03v3 w=1.7u l=0.3u m=1
X2 Y A GND GND nfet_03v3 w=0.85u l=0.3u m=1
X3 Y B GND GND nfet_03v3 w=0.85u l=0.3u m=1
X4 Y C net2 VDD pfet_03v3 w=1.7u l=0.3u m=1
X5 Y C GND GND nfet_03v3 w=0.85u l=0.3u m=1
.ends
.GLOBAL VDD
.GLOBAL GND
