VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp9t3v3__nand3_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__nand3_1 ;
  ORIGIN -5.150 0.000 ;
  SIZE 3.900 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 3.050 6.250 3.350 ;
      LAYER Metal2 ;
        RECT 5.750 3.000 6.250 3.400 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.050 3.050 7.550 3.350 ;
      LAYER Metal2 ;
        RECT 7.050 3.000 7.550 3.400 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 2.210000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 4.400 5.950 5.300 ;
        RECT 7.400 4.450 7.650 5.300 ;
        RECT 7.400 4.400 7.950 4.450 ;
        RECT 5.700 4.150 7.950 4.400 ;
        RECT 6.550 2.700 6.800 4.150 ;
        RECT 5.700 2.450 6.800 2.700 ;
        RECT 5.700 1.050 5.950 2.450 ;
      LAYER Metal2 ;
        RECT 7.450 4.100 7.950 4.500 ;
    END
  END Y
  PIN C
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.500 2.150 8.000 2.450 ;
      LAYER Metal2 ;
        RECT 7.500 2.100 8.000 2.500 ;
    END
  END C
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 5.150 3.150 9.050 6.350 ;
      LAYER Metal1 ;
        RECT 5.150 5.650 9.050 6.350 ;
        RECT 6.550 4.650 6.800 5.650 ;
        RECT 8.250 4.650 8.500 5.650 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 5.150 0.000 9.050 3.150 ;
      LAYER Metal1 ;
        RECT 8.250 0.700 8.500 1.500 ;
        RECT 5.150 0.000 9.050 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.550 1.050 6.800 1.650 ;
        RECT 7.400 1.050 7.650 1.650 ;
  END
END gf180mcu_osu_sc_gp9t3v3__nand3_1
END LIBRARY

