* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__or3_1.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__or3_1 A B C VDD Y VSS
X0 VSS C a_1140_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=17000,540 d=9350,280
X1 VSS A a_1140_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X2 a_1300_720# C a_1140_210# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
**devattr s=34000,880 d=18700,450
X3 a_1140_210# B VSS VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X4 VDD A a_1470_720# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X5 Y a_1140_210# VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=17000,540
X6 a_1470_720# B a_1300_720# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X7 Y a_1140_210# VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=34000,880
.ends

