VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp12t3v3__nor3_1
  CLASS CORE ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__nor3_1 ;
  ORIGIN 0.150 0.000 ;
  SIZE 3.900 BY 8.300 ;
  SYMMETRY XY ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 3.600 0.950 3.900 ;
      LAYER Metal2 ;
        RECT 0.450 3.550 0.950 3.950 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 2.950 1.900 3.250 ;
      LAYER Metal2 ;
        RECT 1.100 2.900 1.600 3.300 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.500 4.250 3.000 4.550 ;
      LAYER Metal2 ;
        RECT 2.500 4.200 3.000 4.600 ;
    END
  END C
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.150 5.100 3.750 8.300 ;
      LAYER Metal1 ;
        RECT -0.150 7.600 3.750 8.300 ;
        RECT 0.400 5.550 0.650 7.600 ;
    END
  END VDD
  PIN Y
    ANTENNADIFFAREA 1.742500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 5.800 2.600 7.250 ;
        RECT 2.000 5.550 2.600 5.800 ;
        RECT 2.000 3.750 2.250 5.550 ;
        RECT 2.000 3.500 2.400 3.750 ;
        RECT 2.150 2.650 2.400 3.500 ;
        RECT 2.150 2.550 3.200 2.650 ;
        RECT 1.250 2.300 3.200 2.550 ;
        RECT 1.250 1.050 1.500 2.300 ;
        RECT 2.500 2.250 3.200 2.300 ;
        RECT 2.950 1.050 3.200 2.250 ;
      LAYER Metal2 ;
        RECT 2.500 2.250 3.000 2.650 ;
    END
  END Y
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 0.700 0.650 1.900 ;
        RECT 2.100 0.700 2.350 1.900 ;
        RECT -0.150 0.000 3.750 0.700 ;
    END
  END VSS
END gf180mcu_osu_sc_gp12t3v3__nor3_1
END LIBRARY

