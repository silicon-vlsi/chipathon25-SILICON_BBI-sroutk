* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__and3_1.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__and3_1 A B Y C VDD VSS
X0 a_250_210# B a_80_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X1 a_n90_210# B VDD VDD pfet_03v3 ad=0.62333p pd=3u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X2 VSS C a_250_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X3 VDD C a_n90_210# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.62333p ps=3u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X4 Y a_n90_210# VSS VSS nfet_03v3 ad=0.4675p pd=2.8u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=18700,560
X5 a_80_210# A a_n90_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.4675p ps=2.8u w=0.85u l=0.3u
**devattr s=18700,560 d=9350,280
X6 Y a_n90_210# VDD VDD pfet_03v3 ad=0.935p pd=4.5u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=37400,900
X7 VDD A a_n90_210# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.62333p ps=3u w=1.7u l=0.3u
**devattr s=37400,900 d=18700,450
C0 a_80_210# a_250_210# 0.05362f
C1 C B 0.09692f
C2 VDD A 0.12462f
C3 a_n90_210# A 0.22916f
C4 VDD B 0.11705f
C5 a_250_210# C 0.02615f
C6 a_n90_210# B 0.18119f
C7 Y C 0.03297f
C8 Y VDD 0.12376f
C9 Y a_n90_210# 0.22425f
C10 a_n90_210# a_80_210# 0.08029f
C11 VDD C 0.08642f
C12 a_n90_210# C 0.14156f
C13 VDD a_n90_210# 0.54827f
C14 B A 0.06819f
C15 Y VSS 0.31925f
C16 C VSS 0.32314f
C17 B VSS 0.28698f
C18 A VSS 0.34197f
C19 VDD VSS 2.13015f
C20 a_250_210# VSS 0.08046f
C21 a_80_210# VSS 0.04401f
C22 a_n90_210# VSS 0.57487f
.ends

