* SPICE3 file created from gf180mcu_osu_sc_gp12t3v3__nand3_1_ext.ext - technology: gf180mcuD

.SUBCKT gf180mcu_osu_sc_gp12t3v3__nand3_1 A B C Y VDD  VSS
X0 VDD A Y VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X1 Y B VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X2 a_250_210# B a_80_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X3 VDD C Y VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X4 VSS C a_250_210# VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X5 a_80_210# A Y VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
C0 Y B 0.13088f
C1 VDD B 0.09252f
C2 VDD Y 0.4416f
C3 B A 0.1103f
C4 Y A 0.2013f
C5 B C 0.09637f
C6 Y C 0.12513f
C7 VDD A 0.1063f
C8 VDD C 0.11076f
C9 VDD VSS 1.79533f
C10 Y VSS 0.56392f 
C11 C VSS 0.61199f 
C12 B VSS 0.51164f 
C13 A VSS 0.57715f 
.ENDS
