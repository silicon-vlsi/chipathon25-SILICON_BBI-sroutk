magic
tech gf180mcuD
timestamp 1755261463
<< nwell >>
rect -17 102 62 166
<< nmos >>
rect 5 21 11 38
rect 22 21 28 38
rect 33 21 39 38
<< pmos >>
rect 2 111 8 145
rect 19 111 25 145
rect 36 111 42 145
<< ndiff >>
rect -8 33 5 38
rect -8 23 -6 33
rect -1 23 5 33
rect -8 21 5 23
rect 11 36 22 38
rect 11 23 14 36
rect 19 23 22 36
rect 11 21 22 23
rect 28 21 33 38
rect 39 36 49 38
rect 39 23 42 36
rect 47 23 49 36
rect 39 21 49 23
<< pdiff >>
rect -8 143 2 145
rect -8 113 -6 143
rect -1 113 2 143
rect -8 111 2 113
rect 8 143 19 145
rect 8 113 11 143
rect 16 113 19 143
rect 8 111 19 113
rect 25 143 36 145
rect 25 113 28 143
rect 33 113 36 143
rect 25 111 36 113
rect 42 143 52 145
rect 42 113 45 143
rect 50 113 52 143
rect 42 111 52 113
<< ndiffc >>
rect -6 23 -1 33
rect 14 23 19 36
rect 42 23 47 36
<< pdiffc >>
rect -6 113 -1 143
rect 11 113 16 143
rect 28 113 33 143
rect 45 113 50 143
<< psubdiff >>
rect 6 12 21 14
rect 6 7 11 12
rect 16 7 21 12
rect 6 5 21 7
rect 30 12 45 14
rect 30 7 35 12
rect 40 7 45 12
rect 30 5 45 7
<< nsubdiff >>
rect 6 159 21 161
rect 6 154 11 159
rect 16 154 21 159
rect 6 152 21 154
rect 30 159 45 161
rect 30 154 35 159
rect 40 154 45 159
rect 30 152 45 154
<< psubdiffcont >>
rect 11 7 16 12
rect 35 7 40 12
<< nsubdiffcont >>
rect 11 154 16 159
rect 35 154 40 159
<< polysilicon >>
rect 2 145 8 150
rect 19 145 25 150
rect 36 145 42 150
rect 2 101 8 111
rect -3 97 8 101
rect -3 61 2 97
rect 19 80 25 111
rect 11 78 25 80
rect 11 72 14 78
rect 20 72 25 78
rect 11 70 25 72
rect -3 59 11 61
rect -3 53 0 59
rect 7 53 11 59
rect -3 50 11 53
rect 5 38 11 50
rect 19 47 25 70
rect 36 67 42 111
rect 36 65 48 67
rect 36 59 40 65
rect 46 59 48 65
rect 36 57 48 59
rect 36 47 42 57
rect 19 43 28 47
rect 22 38 28 43
rect 33 43 42 47
rect 33 38 39 43
rect 5 16 11 21
rect 22 16 28 21
rect 33 16 39 21
<< polycontact >>
rect 14 72 20 78
rect 0 53 7 59
rect 40 59 46 65
<< metal1 >>
rect -17 159 62 166
rect -17 154 11 159
rect 16 154 35 159
rect 40 154 62 159
rect -17 152 62 154
rect -6 143 -1 145
rect -14 108 -1 113
rect 11 143 16 152
rect 11 111 16 113
rect 28 143 33 145
rect -14 91 -9 108
rect 28 91 33 113
rect 45 143 50 152
rect 45 111 50 113
rect -14 85 28 91
rect 34 85 36 91
rect -14 43 -9 85
rect 12 72 14 78
rect 20 72 22 78
rect -2 59 11 61
rect 38 59 40 65
rect 46 59 48 65
rect -2 53 0 59
rect 7 53 11 59
rect -2 51 11 53
rect -14 40 -4 43
rect -14 35 -1 40
rect -6 33 -1 35
rect -6 21 -1 23
rect 14 36 19 38
rect 14 21 19 23
rect 42 36 47 38
rect 42 14 47 23
rect -17 12 62 14
rect -17 7 11 12
rect 16 7 35 12
rect 40 7 62 12
rect -17 0 62 7
<< via1 >>
rect 28 85 34 91
rect 14 72 20 78
rect 40 59 46 65
rect 0 53 7 59
<< metal2 >>
rect 26 91 36 92
rect 26 85 28 91
rect 34 85 36 91
rect 26 84 36 85
rect 12 78 22 79
rect 12 72 14 78
rect 20 72 22 78
rect 12 71 22 72
rect 38 65 48 66
rect -1 59 8 60
rect -1 53 0 59
rect 7 53 8 59
rect 38 59 40 65
rect 46 59 48 65
rect 38 58 48 59
rect -1 52 8 53
<< labels >>
rlabel metal2 17 75 17 75 1 A
port 1 n
rlabel metal2 43 62 43 62 1 B
port 2 n
rlabel via1 31 88 31 88 1 Y
port 3 n
rlabel nsubdiffcont 13 156 13 156 1 VDD
port 4 n
rlabel psubdiffcont 13 9 13 9 1 VSS
port 5 n
flabel metal2 0 59 7 59 5 FreeSans 32 0 0 0 A
flabel metal2 14 78 20 78 5 FreeSans 32 0 0 0 B
flabel metal2 40 65 46 65 5 FreeSans 32 0 0 0 C
flabel metal2 28 91 34 91 5 FreeSans 32 0 0 0 Y
flabel metal1 2 164 36 164 5 FreeSans 32 0 0 0 VDD
flabel metal1 6 3 40 3 1 FreeSans 32 0 0 0 VSS
<< end >>
