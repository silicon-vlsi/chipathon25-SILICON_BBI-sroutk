magic
tech gf180mcuD
timestamp 1755425266
<< nwell >>
rect -17 102 62 166
<< nmos >>
rect 2 21 8 38
rect 19 21 25 38
rect 36 21 42 38
<< pmos >>
rect 2 111 8 145
rect 19 111 25 145
rect 36 111 42 145
<< ndiff >>
rect -8 31 2 38
rect -8 23 -6 31
rect -1 23 2 31
rect -8 21 2 23
rect 8 21 19 38
rect 25 21 36 38
rect 42 36 52 38
rect 42 23 45 36
rect 50 23 52 36
rect 42 21 52 23
<< pdiff >>
rect -8 143 2 145
rect -8 113 -6 143
rect -1 113 2 143
rect -8 111 2 113
rect 8 143 19 145
rect 8 127 11 143
rect 16 127 19 143
rect 8 111 19 127
rect 25 143 36 145
rect 25 113 28 143
rect 33 113 36 143
rect 25 111 36 113
rect 42 143 52 145
rect 42 113 45 143
rect 50 113 52 143
rect 42 111 52 113
<< ndiffc >>
rect -6 23 -1 31
rect 45 23 50 36
<< pdiffc >>
rect -6 113 -1 143
rect 11 127 16 143
rect 28 113 33 143
rect 45 113 50 143
<< psubdiff >>
rect 39 12 52 14
rect 39 7 45 12
rect 50 7 52 12
rect 39 5 52 7
<< nsubdiff >>
rect 6 159 21 161
rect 6 154 11 159
rect 16 154 21 159
rect 6 152 21 154
rect 39 159 52 161
rect 39 154 45 159
rect 50 154 52 159
rect 39 152 52 154
<< psubdiffcont >>
rect 45 7 50 12
<< nsubdiffcont >>
rect 11 154 16 159
rect 45 154 50 159
<< polysilicon >>
rect 2 145 8 150
rect 19 145 25 150
rect 36 145 42 150
rect 2 100 8 111
rect -3 98 8 100
rect -3 92 -1 98
rect 5 92 8 98
rect -3 90 8 92
rect 2 38 8 90
rect 19 52 25 111
rect 14 50 25 52
rect 14 44 16 50
rect 22 44 25 50
rect 14 42 25 44
rect 19 38 25 42
rect 36 80 42 111
rect 36 78 47 80
rect 36 71 39 78
rect 45 71 47 78
rect 36 69 47 71
rect 36 38 42 69
rect 2 16 8 21
rect 19 16 25 21
rect 36 16 42 21
<< polycontact >>
rect -1 92 5 98
rect 16 44 22 50
rect 39 71 45 78
<< metal1 >>
rect -17 159 62 166
rect -17 154 11 159
rect 16 154 45 159
rect 50 154 62 159
rect -17 152 62 154
rect -6 143 -1 145
rect 11 143 16 152
rect 11 125 16 127
rect 28 143 33 145
rect -6 109 -1 113
rect 28 109 33 113
rect 45 143 50 152
rect 45 111 50 113
rect -6 108 33 109
rect -6 107 35 108
rect -6 104 27 107
rect 25 101 27 104
rect 33 101 35 107
rect 25 100 35 101
rect -2 98 6 99
rect -2 92 -1 98
rect 5 92 6 98
rect -2 91 6 92
rect 15 50 23 51
rect 15 44 16 50
rect 22 44 23 50
rect 15 43 23 44
rect 28 33 33 100
rect 38 78 46 79
rect 38 71 39 78
rect 45 71 46 78
rect 38 70 46 71
rect -6 31 33 33
rect -1 28 33 31
rect 45 36 50 38
rect -6 21 -1 23
rect 45 14 50 23
rect -17 12 61 14
rect -17 7 45 12
rect 50 7 61 12
rect -17 0 61 7
<< via1 >>
rect 27 101 33 107
rect -1 92 5 98
rect 16 44 22 50
rect 39 71 45 78
<< metal2 >>
rect 26 107 35 108
rect 26 101 27 107
rect 33 101 35 107
rect 26 100 35 101
rect -2 98 6 99
rect -2 92 -1 98
rect 5 92 6 98
rect -2 91 6 92
rect 38 78 46 79
rect 38 71 39 78
rect 45 71 46 78
rect 38 70 46 71
rect 15 50 23 51
rect 15 44 16 50
rect 22 44 23 50
rect 15 43 23 44
<< labels >>
rlabel nsubdiffcont 13 156 13 156 1 VDD
port 4 n
flabel nwell 2 164 36 164 5 FreeSans 32 0 0 0 VDD
flabel metal1 6 3 40 3 1 FreeSans 32 0 0 0 VSS
rlabel psubdiffcont 47 9 47 9 1 VSS
port 5 n
rlabel nsubdiffcont 47 156 47 156 1 VDD
port 4 n
rlabel metal2 -1 92 5 98 1 A
rlabel via1 27 101 33 107 1 Y
rlabel metal2 39 71 45 78 1 C
rlabel metal2 16 44 22 50 1 B
flabel metal2 21 45 21 49 7 FreeSans 32 0 0 0 B
flabel metal2 40 72 40 77 3 FreeSans 32 0 0 0 C
flabel via1 28 102 32 102 1 FreeSans 32 0 0 0 Y
flabel metal2 0 93 0 97 3 FreeSans 32 0 0 0 A
<< end >>
