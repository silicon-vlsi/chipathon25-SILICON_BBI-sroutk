* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__nor3_1.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__nor3_1 A B C VDD Y VSS
X0 Y A VSS VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=17000,540 d=9350,280
X1 Y C VSS VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=9350,280 d=17000,540
X2 a_1390_720# A VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
**devattr s=34000,880 d=18700,450
X3 VSS B Y VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X4 Y C a_1560_720# VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=34000,880
X5 a_1560_720# B a_1390_720# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
C0 Y C 0.3582f
C1 Y VDD 0.15691f
C2 Y A 0.08406f
C3 Y a_1390_720# 0.0207f
C4 C VDD 0.11629f
C5 A VDD 0.11749f
C6 a_1390_720# VDD 0.01026f
C7 Y B 0.14455f
C8 B C 0.19645f
C9 B VDD 0.08483f
C10 A B 0.06746f
C11 Y a_1560_720# 0.02983f
C12 Y VSS 0.5073f
C13 C VSS 0.33215f
C14 B VSS 0.33068f
C15 A VSS 0.41565f
C16 VDD VSS 1.75173f
.ends

