* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__or3_1.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__or3_1 A B C VDD Y VSS
X0 VSS C a_1140_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=17000,540 d=9350,280
X1 VSS A a_1140_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X2 a_1300_720# C a_1140_210# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
**devattr s=34000,880 d=18700,450
X3 a_1140_210# B VSS VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X4 VDD A a_1470_720# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X5 Y a_1140_210# VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=17000,540
X6 a_1470_720# B a_1300_720# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X7 Y a_1140_210# VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=34000,880
C0 a_1140_210# a_1300_720# 0.11903f
C1 A a_1140_210# 0.14684f
C2 B VDD 0.1132f
C3 a_1470_720# VDD 0.1069f
C4 Y VDD 0.13672f
C5 B a_1140_210# 0.2365f
C6 a_1470_720# a_1140_210# 0.05147f
C7 B C 0.06746f
C8 a_1140_210# Y 0.20607f
C9 a_1140_210# VDD 0.29238f
C10 B A 0.07464f
C11 a_1470_720# a_1300_720# 0.06721f
C12 VDD C 0.12385f
C13 A Y 0.04072f
C14 a_1300_720# VDD 0.0397f
C15 A VDD 0.08867f
C16 a_1140_210# C 0.21649f
C17 Y VSS 0.30794f
C18 A VSS 0.31593f
C19 B VSS 0.28642f
C20 C VSS 0.35179f
C21 VDD VSS 2.1747f
C22 a_1470_720# VSS 0.01192f
C23 a_1300_720# VSS 0.01188f
C24 a_1140_210# VSS 0.82154f
.ends

