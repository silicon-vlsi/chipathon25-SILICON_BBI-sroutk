* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__nor3_1.ext - technology: gf180mcuD

.subckt nor3 A B C VDD Y VSS
X0 Y A VSS VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=17000,540 d=9350,280
X1 Y C VSS VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=9350,280 d=17000,540
X2 a_1390_720# A VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
**devattr s=34000,880 d=18700,450
X3 VSS B Y VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X4 Y C a_1560_720# VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=34000,880
X5 a_1560_720# B a_1390_720# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
.ends

