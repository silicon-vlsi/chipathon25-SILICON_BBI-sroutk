* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__and3_1.ext - technology: gf180mcuD

X0 Y a_9_21# VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X1 VDD C a_9_21# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.595p ps=2.96667u w=1.7u l=0.3u
X2 a_9_21# B VDD VDD pfet_03v3 ad=0.595p pd=2.96667u as=0.4675p ps=2.25u w=1.7u l=0.3u
X3 VDD A a_9_21# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.595p ps=2.96667u w=1.7u l=0.3u
X4 VSS C a_42_21# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X5 a_25_21# A a_9_21# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X6 Y a_9_21# VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X7 a_42_21# B a_25_21# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
C0 A C 0.00152f
C1 B A 0.09405f
C2 Y A 0
C3 C a_9_21# 0.19919f
C4 a_25_21# a_9_21# 0.00723f
C5 a_42_21# a_9_21# 0.00188f
C6 B a_9_21# 0.16365f
C7 Y a_9_21# 0.16617f
C8 A a_9_21# 0.236f
C9 VDD C 0.09443f
C10 B VDD 0.0938f
C11 Y VDD 0.19148f
C12 VDD A 0.10084f
C13 B C 0.11486f
C14 Y C 0.03355f
C15 B a_42_21# 0.00239f
C16 VDD a_9_21# 0.65493f
C17 Y B 0.01334f
C18 a_42_21# VSS 0.00795f
C19 a_25_21# VSS 0.00738f
C20 Y VSS 0.46251f
C21 a_9_21# VSS 1.03872f
C22 C VSS 0.52541f
C23 B VSS 0.51514f
C24 A VSS 0.61257f
C25 VDD VSS 2.09312f
