magic
tech gf180mcuD
magscale 1 5
timestamp 1755251956
<< error_p >>
rect 195 260 245 263
<< nwell >>
rect 0 315 405 635
<< nmos >>
rect 95 105 125 190
rect 180 105 210 190
rect 275 105 305 190
<< pmos >>
rect 110 360 140 530
rect 165 360 195 530
rect 255 360 285 530
<< ndiff >>
rect 45 180 95 190
rect 45 115 55 180
rect 80 115 95 180
rect 45 105 95 115
rect 125 180 180 190
rect 125 115 140 180
rect 165 115 180 180
rect 125 105 180 115
rect 210 180 275 190
rect 210 115 225 180
rect 250 115 275 180
rect 210 105 275 115
rect 305 180 355 190
rect 305 115 320 180
rect 345 115 355 180
rect 305 105 355 115
<< pdiff >>
rect 60 520 110 530
rect 60 370 70 520
rect 95 370 110 520
rect 60 360 110 370
rect 140 360 165 530
rect 195 360 255 530
rect 285 520 345 530
rect 285 370 300 520
rect 325 370 345 520
rect 285 360 345 370
<< ndiffc >>
rect 55 115 80 180
rect 140 115 165 180
rect 225 115 250 180
rect 320 115 345 180
<< pdiffc >>
rect 70 370 95 520
rect 300 370 325 520
<< psubdiff >>
rect 30 60 105 70
rect 30 35 55 60
rect 80 35 105 60
rect 30 25 105 35
rect 150 60 225 70
rect 150 35 175 60
rect 200 35 225 60
rect 150 25 225 35
rect 270 60 345 70
rect 270 35 295 60
rect 320 35 345 60
rect 270 25 345 35
<< nsubdiff >>
rect 30 600 105 610
rect 30 575 55 600
rect 80 575 105 600
rect 30 565 105 575
rect 150 600 225 610
rect 150 575 175 600
rect 200 575 225 600
rect 150 565 225 575
rect 295 600 370 610
rect 295 575 315 600
rect 340 575 370 600
rect 295 565 370 575
<< psubdiffcont >>
rect 55 35 80 60
rect 175 35 200 60
rect 295 35 320 60
<< nsubdiffcont >>
rect 55 575 80 600
rect 175 575 200 600
rect 315 575 340 600
<< polysilicon >>
rect 110 530 140 555
rect 165 530 195 555
rect 255 530 285 555
rect 110 340 140 360
rect 95 315 140 340
rect 165 345 195 360
rect 165 315 210 345
rect 255 340 285 360
rect 255 325 300 340
rect 95 270 125 315
rect 55 260 125 270
rect 55 230 70 260
rect 100 230 125 260
rect 55 220 125 230
rect 95 190 125 220
rect 180 300 210 315
rect 275 315 300 325
rect 275 310 305 315
rect 275 300 345 310
rect 180 290 250 300
rect 180 260 205 290
rect 235 260 250 290
rect 180 250 250 260
rect 275 270 300 300
rect 330 270 345 300
rect 275 260 345 270
rect 180 190 210 250
rect 275 190 305 260
rect 95 80 125 105
rect 180 80 210 105
rect 275 80 305 105
<< polycontact >>
rect 70 230 100 260
rect 205 260 235 290
rect 300 270 330 300
<< metal1 >>
rect 0 600 405 635
rect 0 575 55 600
rect 80 575 175 600
rect 200 575 315 600
rect 340 575 405 600
rect 0 565 405 575
rect 70 520 95 565
rect 70 360 95 370
rect 300 520 325 530
rect 300 350 325 370
rect 300 325 390 350
rect 195 260 205 290
rect 235 260 245 290
rect 290 270 300 300
rect 330 270 340 300
rect 60 230 70 260
rect 100 230 110 260
rect 365 240 390 325
rect 140 215 390 240
rect 55 180 80 190
rect 55 70 80 115
rect 140 180 165 215
rect 140 105 165 115
rect 225 180 250 190
rect 225 70 250 115
rect 320 180 345 215
rect 320 105 345 115
rect 0 60 405 70
rect 0 35 55 60
rect 80 35 175 60
rect 200 35 295 60
rect 320 35 405 60
rect 0 0 405 35
<< via1 >>
rect 205 260 235 290
rect 300 270 330 300
rect 70 230 100 260
<< metal2 >>
rect 290 300 340 305
rect 195 290 245 295
rect 60 260 110 265
rect 60 230 70 260
rect 100 230 110 260
rect 195 260 205 290
rect 235 260 245 290
rect 290 270 300 300
rect 330 270 340 300
rect 290 265 340 270
rect 195 255 245 260
rect 60 225 110 230
<< labels >>
rlabel nsubdiffcont 65 585 65 585 1 VDD
port 4 n
rlabel psubdiffcont 65 45 65 45 1 VSS
port 5 n
rlabel metal2 85 245 85 245 1 A
port 1 n
<< end >>
