magic
tech gf180mcuD
magscale 1 10
timestamp 1755268915
<< error_p >>
rect 1790 480 1810 670
rect 1310 407 1360 410
rect 1310 397 1313 407
rect 1310 363 1313 383
rect 1357 363 1360 407
rect 1310 360 1360 363
rect 779 320 790 331
rect 570 317 620 320
rect 740 317 801 320
rect 570 273 573 317
rect 740 273 743 317
rect 787 309 801 317
rect 787 307 790 309
rect 787 281 790 293
rect 787 273 801 281
rect 570 270 620 273
rect 740 270 801 273
rect 779 259 790 270
rect 830 200 860 220
<< nwell >>
rect 420 342 1910 860
rect 860 340 1910 342
<< pwell >>
rect 420 340 860 342
rect 420 210 1910 340
rect 420 200 480 210
rect 620 200 680 210
rect 710 200 760 210
rect 780 200 1910 210
rect 420 110 1910 200
rect 420 70 480 110
rect 540 70 590 110
rect 620 70 680 110
rect 780 70 1910 110
rect 420 -96 1910 70
rect 860 -100 1910 -96
<< nmos >>
rect 620 110 680 200
<< pmos >>
rect 620 510 680 670
<< mvnmos >>
rect 930 60 1050 220
rect 1160 60 1280 220
rect 1580 60 1700 220
<< mvpmos >>
rect 930 570 1030 670
rect 1160 570 1260 670
rect 1590 480 1690 670
<< ndiff >>
rect 510 180 620 200
rect 510 130 540 180
rect 590 130 620 180
rect 510 110 620 130
rect 680 180 780 200
rect 680 130 710 180
rect 760 130 780 180
rect 680 110 780 130
<< pdiff >>
rect 510 640 620 670
rect 510 590 540 640
rect 590 590 620 640
rect 510 510 620 590
rect 680 640 780 670
rect 680 590 710 640
rect 760 590 780 640
rect 680 510 780 590
<< mvndiff >>
rect 830 190 930 220
rect 830 140 850 190
rect 900 140 930 190
rect 830 60 930 140
rect 1050 190 1160 220
rect 1050 140 1080 190
rect 1130 140 1160 190
rect 1050 60 1160 140
rect 1280 190 1380 220
rect 1280 140 1310 190
rect 1360 140 1380 190
rect 1280 60 1380 140
rect 1470 140 1580 220
rect 1470 90 1500 140
rect 1550 90 1580 140
rect 1470 60 1580 90
rect 1700 190 1810 220
rect 1700 140 1730 190
rect 1780 140 1810 190
rect 1700 60 1810 140
<< mvpdiff >>
rect 830 640 930 670
rect 830 590 850 640
rect 900 590 930 640
rect 830 570 930 590
rect 1030 650 1160 670
rect 1030 600 1070 650
rect 1120 600 1160 650
rect 1030 570 1160 600
rect 1260 640 1380 670
rect 1260 590 1310 640
rect 1360 590 1380 640
rect 1260 570 1380 590
rect 1470 650 1590 670
rect 1470 600 1500 650
rect 1550 600 1590 650
rect 1470 480 1590 600
rect 1690 640 1810 670
rect 1690 590 1730 640
rect 1780 590 1810 640
rect 1690 480 1810 590
<< ndiffc >>
rect 540 130 590 180
rect 710 130 760 180
<< pdiffc >>
rect 540 590 590 640
rect 710 590 760 640
<< mvndiffc >>
rect 850 140 900 190
rect 1080 140 1130 190
rect 1310 140 1360 190
rect 1500 90 1550 140
rect 1730 140 1780 190
<< mvpdiffc >>
rect 850 590 900 640
rect 1070 600 1120 650
rect 1310 590 1360 640
rect 1500 600 1550 650
rect 1730 590 1780 640
<< polysilicon >>
rect 620 670 680 720
rect 930 670 1030 720
rect 1160 670 1260 720
rect 1590 670 1690 720
rect 620 330 680 510
rect 930 480 1030 570
rect 990 410 1030 480
rect 1160 530 1260 570
rect 1160 480 1180 530
rect 1230 480 1260 530
rect 1160 460 1250 480
rect 1300 410 1370 420
rect 990 370 1310 410
rect 1300 360 1310 370
rect 1360 360 1370 410
rect 1590 390 1690 480
rect 1300 350 1370 360
rect 560 320 680 330
rect 560 270 570 320
rect 620 270 680 320
rect 560 260 680 270
rect 730 320 800 330
rect 730 270 740 320
rect 790 280 1050 320
rect 1580 310 1700 390
rect 790 270 800 280
rect 730 260 800 270
rect 620 200 680 260
rect 930 220 1050 280
rect 1160 220 1280 300
rect 1580 260 1610 310
rect 1660 260 1700 310
rect 1580 220 1700 260
rect 620 60 680 110
rect 930 10 1050 60
rect 1160 10 1280 60
rect 1580 10 1700 60
<< polycontact >>
rect 1180 480 1230 530
rect 1310 360 1360 410
rect 570 270 620 320
rect 740 270 790 320
rect 1610 260 1660 310
<< metal1 >>
rect 420 714 1910 834
rect 540 640 590 714
rect 540 520 590 590
rect 710 640 760 660
rect 510 320 650 330
rect 510 270 570 320
rect 620 270 650 320
rect 510 260 650 270
rect 710 320 760 590
rect 850 640 900 660
rect 850 530 900 590
rect 1060 650 1130 714
rect 1060 600 1070 650
rect 1120 600 1130 650
rect 1060 580 1130 600
rect 1310 640 1360 660
rect 850 480 1180 530
rect 1230 480 1260 530
rect 710 270 740 320
rect 540 180 590 200
rect 540 50 590 130
rect 710 180 760 270
rect 710 110 760 130
rect 850 190 900 480
rect 1310 410 1360 590
rect 1490 650 1560 714
rect 1490 600 1500 650
rect 1550 600 1560 650
rect 1490 580 1560 600
rect 1730 640 1780 660
rect 1310 320 1360 360
rect 1310 310 1680 320
rect 1310 260 1610 310
rect 1660 260 1680 310
rect 1310 250 1680 260
rect 850 110 900 140
rect 1080 190 1130 220
rect 1080 50 1130 140
rect 1310 190 1360 250
rect 1730 190 1780 590
rect 1310 110 1360 140
rect 1500 140 1550 160
rect 1730 100 1780 140
rect 1500 50 1550 90
rect 420 -70 1910 50
<< labels >>
rlabel metal1 1730 350 1780 400 1 Y
rlabel polycontact 570 270 620 320 1 A
<< properties >>
string FIXED_BBOX -10 -10 774 774
<< end >>
