* SPICE3 file created from gf180mcu_osu_sc_gp12t3v3__nor3_1_lay.ext - technology: gf180mcuD

X0 a_220_210# a_60_700# VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X1 VSS a_270_570# a_220_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X2 a_330_1110# a_270_570# a_220_1110# VDD pfet_03v3 ad=0.2125p pd=1.95u as=0.2125p ps=1.95u w=1.7u l=0.3u
X3 a_220_210# a_380_1020# VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X4 a_220_210# a_380_1020# a_330_1110# VDD pfet_03v3 ad=1.105p pd=4.7u as=0.2125p ps=1.95u w=1.7u l=0.3u
X5 a_220_1110# a_60_700# VDD VDD pfet_03v3 ad=0.2125p pd=1.95u as=0.85p ps=4.4u w=1.7u l=0.3u
