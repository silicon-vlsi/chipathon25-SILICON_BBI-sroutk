* SPICE3 file created from gf180mcu_osu_sc_gp12t3v3__nor3_1_ext_lvs.ext - technology: gf180mcuD

X0 net3 A VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X1 VSS B net3 VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X2 a_330_1110# B a_220_1110# VDD pfet_03v3 ad=0.2125p pd=1.95u as=0.2125p ps=1.95u w=1.7u l=0.3u
X3 net3 C VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X4 net3 C a_330_1110# VDD pfet_03v3 ad=0.85p pd=4.4u as=0.2125p ps=1.95u w=1.7u l=0.3u
X5 a_220_1110# A VDD VDD pfet_03v3 ad=0.2125p pd=1.95u as=0.85p ps=4.4u w=1.7u l=0.3u
