* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__nor3_1.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp12t3v3__nor3_1 A B C VDD Y VSS
X0 Y A VSS VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=17000,540 d=9350,280
X1 VSS B Y VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X2 a_330_1110# B a_220_1110# VDD pfet_03v3 ad=0.2125p pd=1.95u as=0.2125p ps=1.95u w=1.7u l=0.3u
**devattr s=8500,390 d=8500,390
X3 Y C VSS VSS nfet_03v3 ad=0.2975p pd=1.83333u as=0.2975p ps=1.83333u w=0.85u l=0.3u
**devattr s=9350,280 d=17000,540
X4 Y C a_330_1110# VDD pfet_03v3 ad=0.85p pd=4.4u as=0.2125p ps=1.95u w=1.7u l=0.3u
**devattr s=8500,390 d=34000,880
X5 a_220_1110# A VDD VDD pfet_03v3 ad=0.2125p pd=1.95u as=0.85p ps=4.4u w=1.7u l=0.3u
**devattr s=34000,880 d=8500,390
C0 A B 0.19808f
C1 VDD Y 0.11209f
C2 C Y 0.19895f
C3 VDD C 0.14998f
C4 A Y 0.03661f
C5 A VDD 0.1056f
C6 Y B 0.20803f
C7 VDD B 0.08275f
C8 C B 0.10302f
C9 Y VSS 0.79765f
C10 C VSS 0.62466f
C11 B VSS 0.52627f
C12 A VSS 0.60905f
C13 VDD VSS 1.80377f
.ends

