* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__and3_1.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp12t3v3__and3_1 A B Y C VDD VSS
X0 VDD A a_90_210# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.595p ps=2.96667u w=1.7u l=0.3u
**devattr s=34000,880 d=18700,450
X1 Y a_90_210# VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=34000,880
X2 a_250_210# A a_90_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
**devattr s=17000,540 d=9350,280
X3 a_90_210# B VDD VDD pfet_03v3 ad=0.595p pd=2.96667u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X4 a_420_210# B a_250_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X5 VSS C a_420_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X6 Y a_90_210# VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=17000,540
X7 VDD C a_90_210# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.595p ps=2.96667u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
C0 B Y 0.01334f
C1 a_90_210# Y 0.16617f
C2 B A 0.09405f
C3 A a_90_210# 0.236f
C4 VDD C 0.09443f
C5 B VDD 0.0938f
C6 B C 0.11486f
C7 VDD a_90_210# 0.65493f
C8 C a_90_210# 0.19919f
C9 VDD Y 0.19148f
C10 C Y 0.03355f
C11 VDD A 0.10084f
C12 B a_90_210# 0.16365f
C13 Y VSS 0.46251f
C14 C VSS 0.52541f
C15 B VSS 0.51514f
C16 A VSS 0.61257f
C17 VDD VSS 2.09312f
C18 a_90_210# VSS 1.03872f
.ends

