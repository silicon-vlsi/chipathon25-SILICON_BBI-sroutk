VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp12t3v3__nor3_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__nor3_1 ;
  ORIGIN 0.150 0.000 ;
  SIZE 3.900 BY 8.300 ;
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.150 5.100 3.750 8.300 ;
      LAYER Metal1 ;
        RECT -0.150 7.600 3.750 8.300 ;
        RECT 0.400 5.550 0.650 7.600 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 0.700 0.650 1.900 ;
        RECT 2.100 0.700 2.350 1.900 ;
        RECT -0.150 0.000 3.750 0.700 ;
    END
  END VSS
  PIN Y
    ANTENNADIFFAREA 1.742500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 5.400 2.600 7.250 ;
        RECT 2.200 5.150 2.600 5.400 ;
        RECT 2.200 2.600 2.450 5.150 ;
        RECT 2.900 2.650 3.250 2.700 ;
        RECT 2.800 2.600 3.300 2.650 ;
        RECT 2.200 2.550 3.300 2.600 ;
        RECT 1.250 2.300 3.300 2.550 ;
        RECT 1.250 1.050 1.500 2.300 ;
        RECT 2.800 2.250 3.300 2.300 ;
        RECT 2.950 1.050 3.200 2.250 ;
      LAYER Metal2 ;
        RECT 2.800 2.250 3.300 2.650 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 2.800 4.100 3.300 4.400 ;
        RECT 0.300 3.600 0.800 3.900 ;
        RECT 1.400 2.950 1.900 3.250 ;
      LAYER Metal2 ;
        RECT 2.800 4.050 3.300 4.450 ;
        RECT 0.300 3.550 0.800 3.950 ;
        RECT 1.400 2.900 1.900 3.300 ;
  END
END gf180mcu_osu_sc_gp12t3v3__nor3_1
END LIBRARY

