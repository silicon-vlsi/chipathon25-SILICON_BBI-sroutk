** sch_path: /foss/designs/work/xschem/gf180mcu_osu_sc_gp12t3v3__nor3_1.sch
.subckt gf180mcu_osu_sc_gp12t3v3__nor3_1 A B C VDD VSS Y VSS VSS
*.PININFO A:I B:I C:I VDD:B VSS:B Y:O VSS:B VSS:B
X1 net2 A VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X2 net1 B net2 VDD pfet_03v3 w=1.7u l=0.3u m=1
X3 Y C net1 VDD pfet_03v3 w=1.7u l=0.3u m=1
X4 Y A VSS VSS nfet_03v3 w=0.85u l=0.3u m=1
X5 Y B VSS VSS nfet_03v3 w=0.85u l=0.3u m=1
X6 Y C VSS VSS nfet_03v3 w=0.85u l=0.3u m=1
.ends
