** sch_path: /foss/designs/work/xschem/TB_nand1_3.sch
**.subckt TB_nand1_3

.PARAM PAR_CLOAD=5f
.PARAM PAR_SLEW=100p
.PARAM PAR_PERIOD=10n
.PARAM PAR_TSTOP=PAR_PERIOD

.INCLUDE ../../core_digital/gf180mcu_osu_sc_gp12t3v3/cells/nand3/gf180mcu_osu_sc_gp12t3v3__nand3_1.spice

**netlist
Xnand 	A B Y C VDD VSS gf180mcu_osu_sc_gp12t3v3__nand3_1
Cload   Y     	VSS   50f

**Sources
Vdc   	VDD   	VSS   	3.3
VinA   	A    	VSS   	0 	PULSE(0 3.3 1n 1p 1p 5n 10n)
VinB   	B    	VSS   	0	PULSE(0 3.3 2n 1p 1p 5n 10n)
VinC   	C    	VSS   	0	PULSE(0 3.3 3n 1p 1p 5n 10n)
Vgnd	

** Rise/Fall 10-90%
.MEASURE TRAN tr1090 TRIG v(Y) VAL='0.1*1.8' RISE=1 TARG v(Y) VAL='0.9*1.8' RISE=1
.MEASURE TRAN tf9010 TRIG v(Y) VAL='0.9*1.8' FALL=1 TARG v(Y) VAL='0.1*1.8' FALL=1

** Delay Rise Fall
.MEASURE TRAN tdrise TRIG v(A)  VAL='0.5*1.8' RISE=1 TARG v(Y) VAL='0.5*1.8' RISE=1
.MEASURE TRAN tdfall TRIG v(A)  VAL='0.5*1.8' FALL=1 TARG v(Y) VAL='0.5*1.8' FALL=1

.control
save all
op
tran 1p 20n
.endc



.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends
.end
