magic
tech gf180mcuD
timestamp 1755549038
<< nwell >>
rect -10 63 81 127
<< nmos >>
rect 12 21 18 38
rect 29 21 35 38
rect 51 21 57 38
<< pmos >>
rect 12 72 18 106
rect 29 72 35 106
rect 51 72 57 106
<< ndiff >>
rect -1 36 12 38
rect -1 23 1 36
rect 6 23 12 36
rect -1 21 12 23
rect 18 36 29 38
rect 18 23 21 36
rect 26 23 29 36
rect 18 21 29 23
rect 35 36 51 38
rect 35 23 40 36
rect 45 23 51 36
rect 35 21 51 23
rect 57 36 71 38
rect 57 23 64 36
rect 69 23 71 36
rect 57 21 71 23
<< pdiff >>
rect 2 104 12 106
rect 2 74 4 104
rect 9 74 12 104
rect 2 72 12 74
rect 18 72 29 106
rect 35 72 51 106
rect 57 104 69 106
rect 57 80 62 104
rect 67 80 69 104
rect 57 72 69 80
<< ndiffc >>
rect 1 23 6 36
rect 21 23 26 36
rect 40 23 45 36
rect 64 23 69 36
<< pdiffc >>
rect 4 74 9 104
rect 62 80 67 104
<< psubdiff >>
rect -5 12 10 14
rect -5 7 0 12
rect 5 7 10 12
rect -5 5 10 7
rect 35 12 50 14
rect 35 7 40 12
rect 45 7 50 12
rect 35 5 50 7
rect 61 12 76 14
rect 61 7 66 12
rect 71 7 76 12
rect 61 5 76 7
<< nsubdiff >>
rect 6 120 21 122
rect 6 115 11 120
rect 16 115 21 120
rect 6 113 21 115
rect 30 120 45 122
rect 30 115 35 120
rect 40 115 45 120
rect 30 113 45 115
rect 59 120 74 122
rect 59 115 63 120
rect 68 115 74 120
rect 59 113 74 115
<< psubdiffcont >>
rect 0 7 5 12
rect 40 7 45 12
rect 66 7 71 12
<< nsubdiffcont >>
rect 11 115 16 120
rect 35 115 40 120
rect 63 115 68 120
<< polysilicon >>
rect 12 106 18 111
rect 29 106 35 111
rect 51 106 57 111
rect 12 60 18 72
rect 4 58 18 60
rect 4 52 7 58
rect 13 52 18 58
rect 4 50 18 52
rect 12 38 18 50
rect 29 54 35 72
rect 51 62 57 72
rect 51 60 65 62
rect 51 54 56 60
rect 62 54 65 60
rect 29 52 43 54
rect 29 46 34 52
rect 40 46 43 52
rect 29 44 43 46
rect 51 52 65 54
rect 29 38 35 44
rect 51 38 57 52
rect 12 16 18 21
rect 29 16 35 21
rect 51 16 57 21
<< polycontact >>
rect 7 52 13 58
rect 56 54 62 60
rect 34 46 40 52
<< metal1 >>
rect -10 120 81 127
rect -10 115 11 120
rect 16 115 35 120
rect 40 115 63 120
rect 68 115 81 120
rect -10 113 81 115
rect 4 104 9 113
rect 4 72 9 74
rect 62 104 67 106
rect 62 74 67 80
rect 62 71 66 74
rect 21 68 66 71
rect 72 68 74 74
rect 21 66 67 68
rect 5 52 7 58
rect 13 52 15 58
rect 1 36 6 38
rect 1 14 6 23
rect 21 36 26 66
rect 54 54 56 60
rect 62 54 64 60
rect 32 46 34 52
rect 40 46 42 52
rect 21 21 26 23
rect 40 36 45 38
rect 40 14 45 23
rect 64 36 69 38
rect 64 21 69 23
rect -10 12 81 14
rect -10 7 0 12
rect 5 7 40 12
rect 45 7 66 12
rect 71 7 81 12
rect -10 0 81 7
<< via1 >>
rect 66 68 72 74
rect 7 52 13 58
rect 56 54 62 60
rect 34 46 40 52
<< metal2 >>
rect 64 74 74 75
rect 64 68 66 74
rect 72 68 74 74
rect 64 67 74 68
rect 54 60 64 61
rect 5 58 15 59
rect 5 52 7 58
rect 13 52 15 58
rect 54 54 56 60
rect 62 54 64 60
rect 54 53 64 54
rect 5 51 15 52
rect 32 52 42 53
rect 32 46 34 52
rect 40 46 42 52
rect 32 45 42 46
<< labels >>
rlabel nsubdiffcont 13 117 13 117 1 VDD
port 4 n
<< end >>
