VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp9t3v3__ant
  CLASS CORE ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__ant ;
  ORIGIN -2.550 0.000 ;
  SIZE 1.750 BY 6.350 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN Y1
    ANTENNADIFFAREA 0.637500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.300 2.800 3.550 5.300 ;
        RECT 3.200 2.400 3.600 2.800 ;
        RECT 3.300 1.050 3.550 2.400 ;
      LAYER Metal2 ;
        RECT 3.200 2.400 3.600 2.800 ;
    END
  END Y1
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 2.550 3.150 4.300 6.350 ;
      LAYER Metal1 ;
        RECT 2.550 5.650 4.300 6.350 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.550 0.000 4.300 0.700 ;
    END
  END VSS
END gf180mcu_osu_sc_gp9t3v3__ant
END LIBRARY

