VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp9t3v3__or3_1
  CLASS CORE ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__or3_1 ;
  ORIGIN -5.250 0.000 ;
  SIZE 5.000 BY 6.350 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.800 2.400 8.300 2.700 ;
      LAYER Metal2 ;
        RECT 7.800 2.350 8.300 2.750 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.150 3.100 7.650 3.400 ;
      LAYER Metal2 ;
        RECT 7.150 3.050 7.650 3.450 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 3.100 6.350 3.400 ;
      LAYER Metal2 ;
        RECT 5.850 3.050 6.350 3.450 ;
    END
  END C
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 5.250 3.150 10.250 6.350 ;
      LAYER Metal1 ;
        RECT 5.250 5.650 10.250 6.350 ;
        RECT 8.350 4.400 8.600 5.650 ;
    END
  END VDD
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.200 2.700 9.450 5.300 ;
        RECT 9.100 2.400 9.600 2.700 ;
        RECT 9.200 1.050 9.450 2.400 ;
      LAYER Metal2 ;
        RECT 9.100 2.350 9.600 2.750 ;
    END
  END Y
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.650 0.700 6.900 1.550 ;
        RECT 8.350 0.700 8.600 1.550 ;
        RECT 5.250 0.000 10.250 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 5.800 4.050 6.050 5.300 ;
        RECT 6.650 4.400 6.900 5.300 ;
        RECT 7.500 4.400 7.750 5.300 ;
        RECT 5.800 3.800 8.850 4.050 ;
        RECT 6.650 2.050 6.900 3.800 ;
        RECT 8.550 3.000 8.850 3.800 ;
        RECT 5.800 1.800 7.750 2.050 ;
        RECT 5.800 1.050 6.050 1.800 ;
        RECT 7.500 1.050 7.750 1.800 ;
  END
END gf180mcu_osu_sc_gp9t3v3__or3_1
END LIBRARY

