** sch_path: /foss/designs/works/xschem/TB_3input_nor.sch
**.subckt TB_3input_nor
**** begin user architecture code


.INCLUDE 3input_nor.spice
**Netlist
Xnor A B C VDD VSS Y VSS VSS 3input_nor
Cload Y VSS 50f

**Sources
VDD VDD VSS 3.3
VSS VSS 0 0
VinA A VSS PULSE(0 3.3 0 1p 1p 10n 20n)
VinB B VSS PULSE(0 3.3 2n 1p 1p 20n 40n)
VinC C VSS PULSE(0 3.3 4n 1p 1p 40n 80n)


.param VDD=3.3

* Output rise/fall (10-90% and 90-10%)
.MEASURE TRAN tr1090_Y  TRIG v(Y) VAL='0.1*VDD'  RISE=1 TARG v(Y) VAL='0.9*VDD' RISE=1
.MEASURE TRAN tf9010_Y  TRIG v(Y) VAL='0.9*VDD'  FALL=1 TARG v(Y) VAL='0.1*VDD' FALL=1

* Propagation delays A -> Y

.MEASURE TRAN tdrise_A TRIG v(A) VAL='0.5*VDD' FALL=1 TARG v(Y) VAL='0.5*VDD' RISE=1

.MEASURE TRAN tdfall_A TRIG v(A) VAL='0.5*VDD' RISE=1 TARG v(Y) VAL='0.5*VDD' FALL=1

* Propagation delays B -> Y

.MEASURE TRAN tdrise_B TRIG v(B) VAL='0.5*VDD' FALL=1 TARG v(Y) VAL='0.5*VDD' RISE=1
.MEASURE TRAN tdfall_B TRIG v(B) VAL='0.5*VDD' RISE=1 TARG v(Y) VAL='0.5*VDD' FALL=1

* Propagation delays C -> Y
.MEASURE TRAN tdrise_C TRIG v(C) VAL='0.5*VDD' FALL=1 TARG v(Y) VAL='0.5*VDD' RISE=1
.MEASURE TRAN tdfall_C TRIG v(C) VAL='0.5*VDD' RISE=1 TARG v(Y) VAL='0.5*VDD' FALL=1



.control
save all
op
tran 0.5n 160n
plot v(A) v(B) v(C) v(Y)
*write test_nfet_03v3.raw
.endc
.end



.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends
.end
