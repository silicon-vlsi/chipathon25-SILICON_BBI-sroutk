* SPICE3 file created from gf180mcu_osu_sc_gp12t3v3__nor3_1_ext.ext - technology: gf180mcuD

X0 net3 A VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X1 VSS B net3 VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X2 a_330_1110# B a_220_1110# VDD pfet_03v3 ad=0.2125p pd=1.95u as=0.2125p ps=1.95u w=1.7u l=0.3u
X3 net3 C VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X4 net3 C a_330_1110# VDD pfet_03v3 ad=0.85p pd=4.4u as=0.2125p ps=1.95u w=1.7u l=0.3u
X5 a_220_1110# A VDD VDD pfet_03v3 ad=0.2125p pd=1.95u as=0.85p ps=4.4u w=1.7u l=0.3u
C0 net3 C 0.1677f
C1 A VDD 0.11248f
C2 A B 0.19643f
C3 A net3 0.03072f
C4 VDD B 0.07962f
C5 net3 VDD 0.10733f
C6 VDD C 0.16048f
C7 net3 B 0.17299f
C8 B C 0.10301f
C9 VDD VSS 1.80192f
C10 net3 VSS 0.80093f **FLOATING
C11 C VSS 0.67281f **FLOATING
C12 B VSS 0.50587f **FLOATING
C13 A VSS 0.6389f **FLOATING
