magic
tech gf180mcuD
timestamp 1757661304
<< nwell >>
rect -17 83 61 166
<< nmos >>
rect 2 21 8 38
rect 19 21 25 38
rect 36 21 42 38
<< pmos >>
rect 2 111 8 145
rect 19 111 25 145
rect 36 111 42 145
<< ndiff >>
rect -8 28 2 38
rect -8 23 -6 28
rect -1 23 2 28
rect -8 21 2 23
rect 8 21 19 38
rect 25 21 36 38
rect 42 36 52 38
rect 42 23 45 36
rect 50 23 52 36
rect 42 21 52 23
<< pdiff >>
rect -8 143 2 145
rect -8 113 -6 143
rect -1 113 2 143
rect -8 111 2 113
rect 8 143 19 145
rect 8 127 11 143
rect 16 127 19 143
rect 8 111 19 127
rect 25 143 36 145
rect 25 113 28 143
rect 33 113 36 143
rect 25 111 36 113
rect 42 143 52 145
rect 42 113 45 143
rect 50 113 52 143
rect 42 111 52 113
<< ndiffc >>
rect -6 23 -1 28
rect 45 23 50 36
<< pdiffc >>
rect -6 113 -1 143
rect 11 127 16 143
rect 28 113 33 143
rect 45 113 50 143
<< psubdiff >>
rect 38 12 53 14
rect 38 7 43 12
rect 48 7 53 12
rect 38 5 53 7
<< nsubdiff >>
rect 6 159 21 161
rect 6 154 11 159
rect 16 154 21 159
rect 6 152 21 154
rect 38 159 53 161
rect 38 154 43 159
rect 48 154 53 159
rect 38 152 53 154
<< psubdiffcont >>
rect 43 7 48 12
<< nsubdiffcont >>
rect 11 154 16 159
rect 43 154 48 159
<< polysilicon >>
rect 2 145 8 150
rect 19 145 25 150
rect 36 145 42 150
rect 2 100 8 111
rect -3 98 8 100
rect -3 92 -1 98
rect 5 92 8 98
rect -3 90 8 92
rect 2 38 8 90
rect 19 58 25 111
rect 14 56 25 58
rect 14 50 16 56
rect 22 50 25 56
rect 14 48 25 50
rect 19 38 25 48
rect 36 82 42 111
rect 36 80 49 82
rect 36 74 41 80
rect 47 74 49 80
rect 36 72 49 74
rect 36 38 42 72
rect 2 16 8 21
rect 19 16 25 21
rect 36 16 42 21
<< polycontact >>
rect -1 92 5 98
rect 16 50 22 56
rect 41 74 47 80
<< metal1 >>
rect -17 159 61 166
rect -17 154 11 159
rect 16 154 43 159
rect 48 154 61 159
rect -17 152 61 154
rect -6 143 -1 145
rect 11 143 16 152
rect 11 125 16 127
rect 28 143 33 145
rect -6 109 -1 113
rect 28 109 33 113
rect 45 143 50 152
rect 45 111 50 113
rect -6 108 35 109
rect -6 104 27 108
rect 25 102 27 104
rect 33 102 35 108
rect 25 100 35 102
rect -2 98 6 99
rect -2 92 -1 98
rect 5 92 6 98
rect -2 91 6 92
rect 28 70 33 100
rect 40 80 48 81
rect 40 74 41 80
rect 47 74 48 80
rect 40 73 48 74
rect -6 65 33 70
rect -6 28 -1 65
rect 12 56 20 57
rect 12 50 13 56
rect 22 50 24 56
rect 12 49 20 50
rect -6 21 -1 23
rect 45 36 50 38
rect 45 14 50 23
rect -17 12 61 14
rect -17 7 43 12
rect 48 7 61 12
rect -17 0 61 7
<< via1 >>
rect 27 102 33 108
rect -1 92 5 98
rect 41 74 47 80
rect 13 50 16 56
rect 16 50 19 56
<< metal2 >>
rect 26 108 34 109
rect 26 102 27 108
rect 33 102 34 108
rect 26 101 34 102
rect -2 98 6 99
rect -2 92 -1 98
rect 5 92 6 98
rect -2 91 6 92
rect 40 80 48 81
rect 40 74 41 80
rect 47 74 48 80
rect 40 73 48 74
rect 12 56 20 57
rect 12 50 13 56
rect 19 50 20 56
rect 12 49 20 50
<< labels >>
flabel metal2 -2 91 6 99 0 FreeSans 48 0 0 0 A
port 1 nsew
flabel metal1 -6 155 6 162 0 FreeSans 48 0 0 0 VDD
port 5 nsew
flabel metal1 -6 4 6 11 0 FreeSans 48 0 0 0 VSS
port 6 nsew
flabel metal2 12 49 20 57 0 FreeSans 48 0 0 0 B
port 2 nsew
flabel metal2 26 101 34 109 0 FreeSans 48 0 0 0 Y
port 3 nsew
flabel metal2 40 73 48 81 0 FreeSans 48 0 0 0 C
port 4 nsew
<< properties >>
string FIXED_BBOX -17 0 61 166
<< end >>
