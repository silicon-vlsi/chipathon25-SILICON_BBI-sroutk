VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp9t3v3__nor3_1
  CLASS CORE ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__nor3_1 ;
  ORIGIN -5.700 0.000 ;
  SIZE 3.900 BY 6.350 ;
  SYMMETRY XY ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.300 2.150 6.800 2.450 ;
      LAYER Metal2 ;
        RECT 6.300 2.100 6.800 2.500 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 2.150 8.100 2.450 ;
      LAYER Metal2 ;
        RECT 7.600 2.100 8.100 2.500 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.200 3.400 8.500 3.450 ;
        RECT 7.650 3.100 8.550 3.400 ;
        RECT 7.650 3.050 8.500 3.100 ;
        RECT 7.650 2.800 8.050 3.050 ;
      LAYER Metal2 ;
        RECT 7.650 2.800 8.050 3.200 ;
    END
  END C
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 5.700 3.150 9.600 6.350 ;
      LAYER Metal1 ;
        RECT 5.700 5.650 9.600 6.350 ;
        RECT 6.250 4.450 6.500 5.650 ;
    END
  END VDD
  PIN Y
    ANTENNADIFFAREA 1.742500 ;
    PORT
      LAYER Metal1 ;
        RECT 7.650 4.150 8.050 4.500 ;
        RECT 8.800 4.150 9.050 5.300 ;
        RECT 7.100 3.900 9.050 4.150 ;
        RECT 7.100 1.050 7.350 3.900 ;
        RECT 8.800 1.050 9.050 3.900 ;
      LAYER Metal2 ;
        RECT 7.650 4.100 8.050 4.500 ;
    END
  END Y
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.250 0.700 6.500 1.500 ;
        RECT 7.950 0.700 8.200 1.500 ;
        RECT 5.700 0.000 9.600 0.700 ;
    END
  END VSS
END gf180mcu_osu_sc_gp9t3v3__nor3_1
END LIBRARY

