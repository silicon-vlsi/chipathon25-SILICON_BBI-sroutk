VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp9t3v3__and3_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__and3_1 ;
  ORIGIN 0.900 0.000 ;
  SIZE 4.900 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT -0.200 3.100 0.300 3.400 ;
      LAYER Metal2 ;
        RECT -0.200 3.050 0.300 3.450 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.050 3.100 1.550 3.400 ;
      LAYER Metal2 ;
        RECT 1.050 3.050 1.550 3.450 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.100 2.450 3.350 5.300 ;
        RECT 3.100 2.150 3.700 2.450 ;
        RECT 3.100 1.050 3.350 2.150 ;
      LAYER Metal2 ;
        RECT 3.150 2.100 3.650 2.500 ;
    END
  END Y
  PIN C
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 2.150 2.000 2.450 ;
      LAYER Metal2 ;
        RECT 1.500 2.100 2.000 2.500 ;
    END
  END C
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.900 3.150 4.000 6.350 ;
      LAYER Metal1 ;
        RECT -0.900 5.650 4.000 6.350 ;
        RECT 0.550 4.600 0.800 5.650 ;
        RECT 2.250 4.600 2.500 5.650 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 0.700 2.500 1.500 ;
        RECT -0.900 0.000 3.950 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT -0.300 4.200 -0.050 5.300 ;
        RECT 1.400 4.200 1.650 5.300 ;
        RECT -0.300 3.950 2.750 4.200 ;
        RECT 0.550 2.500 0.800 3.950 ;
        RECT 2.450 3.000 2.750 3.950 ;
        RECT -0.300 2.250 0.800 2.500 ;
        RECT -0.300 1.050 -0.050 2.250 ;
        RECT 0.550 1.050 0.800 1.750 ;
        RECT 1.400 1.050 1.650 1.750 ;
  END
END gf180mcu_osu_sc_gp9t3v3__and3_1
END LIBRARY

