* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__and3_2.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__and3_2 A B Y C VDD VSS
X0 VDD a_n90_210# Y VDD pfet_03v3 ad=0.561p pd=2.7u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=37400,900
X1 a_250_210# B a_80_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X2 a_n90_210# B VDD VDD pfet_03v3 ad=0.62333p pd=3u as=0.561p ps=2.7u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X3 VSS C a_250_210# VSS nfet_03v3 ad=0.31167p pd=1.86667u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X4 VDD C a_n90_210# VDD pfet_03v3 ad=0.561p pd=2.7u as=0.62333p ps=3u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X5 Y a_n90_210# VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.31167p ps=1.86667u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X6 a_80_210# A a_n90_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.4675p ps=2.8u w=0.85u l=0.3u
**devattr s=18700,560 d=9350,280
X7 Y a_n90_210# VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.561p ps=2.7u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X8 VSS a_n90_210# Y VSS nfet_03v3 ad=0.31167p pd=1.86667u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=18700,560
X9 VDD A a_n90_210# VDD pfet_03v3 ad=0.561p pd=2.7u as=0.62333p ps=3u w=1.7u l=0.3u
**devattr s=37400,900 d=18700,450
C0 VDD C 0.0892f
C1 a_n90_210# a_80_210# 0.08029f
C2 VDD A 0.12462f
C3 a_n90_210# VDD 0.66454f
C4 a_250_210# B 0.01256f
C5 B C 0.07434f
C6 Y C 0.03883f
C7 B A 0.06768f
C8 a_n90_210# B 0.2086f
C9 Y a_n90_210# 0.32644f
C10 B VDD 0.11841f
C11 a_n90_210# C 0.13849f
C12 Y VDD 0.19103f
C13 a_80_210# a_250_210# 0.05362f
C14 a_n90_210# A 0.22916f
C15 Y VSS 0.32384f
C16 C VSS 0.30028f
C17 B VSS 0.28997f
C18 A VSS 0.34197f
C19 VDD VSS 2.48934f
C20 a_250_210# VSS 0.08232f
C21 a_80_210# VSS 0.04401f
C22 a_n90_210# VSS 0.83314f
.ends

