* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__and3_1.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp12t3v3__and3_1 A B Y C VDD VSS
X0 VDD A a_90_210# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.595p ps=2.96667u w=1.7u l=0.3u
**devattr s=34000,880 d=18700,450
X1 Y a_90_210# VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=34000,880
X2 a_250_210# A a_90_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
**devattr s=17000,540 d=9350,280
X3 a_90_210# B VDD VDD pfet_03v3 ad=0.595p pd=2.96667u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X4 a_420_210# B a_250_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X5 VSS C a_420_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X6 Y a_90_210# VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=17000,540
X7 VDD C a_90_210# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.595p ps=2.96667u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
C0 Y C 0.03304f
C1 VDD a_90_210# 0.64996f
C2 B C 0.11628f
C3 C a_90_210# 0.19229f
C4 A B 0.09405f
C5 A a_90_210# 0.24626f
C6 Y B 0.01334f
C7 Y a_90_210# 0.31514f
C8 VDD C 0.09833f
C9 A VDD 0.10605f
C10 Y VDD 0.2214f
C11 B a_90_210# 0.16524f
C12 VDD B 0.09846f
C13 Y VSS 0.45963f
C14 C VSS 0.50452f
C15 B VSS 0.50956f
C16 A VSS 0.60717f
C17 VDD VSS 2.14325f
C18 a_90_210# VSS 1.0252f
.ends

