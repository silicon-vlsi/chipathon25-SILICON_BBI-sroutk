** sch_path: /foss/designs/work/xschem/tb_gf180mcu_osu_sc_gp9t3v3__and3_2.sch
**.subckt tb_gf180mcu_osu_sc_gp9t3v3__and3_2
**** begin user architecture code



.INCLUDE gf180mcu_osu_sc_gp9t3v3__and3_2.spice

**Netlist
Xand A B Y C gf180mcu_osu_sc_gp9t3v3__and3_2
Cload 	Y	GND	50F

.PARAM VDD=3.3

**Sources
Vdc	VDD	GND	3.3
VinA	A 	GND	0	PULSE(0 3.3 0 1p 1p 5n 10n)
VinB	B 	GND	0	PULSE(0 3.3 2n 1p 1p 20n 40n)
VinC	C 	GND	0	PULSE(0 3.3 4n 1p 1p 50n 100n)

** Rise/Fall 10-90%
.MEASURE TRAN tr1090 TRIG v(Y) VAL='0.1*VDD' RISE=1 TARG v(Y) VAL='0.9*VDD' RISE=1
.MEASURE TRAN tf9010 TRIG v(Y) VAL='0.9*VDD' FALL=1 TARG v(Y) VAL='0.1*VDD' FALL=1

** Delay Rise Fall
.MEASURE TRAN tdriseA TRIG v(A)  VAL='0.5*VDD' RISE=1 TARG v(Y) VAL='0.5*VDD' RISE=1
.MEASURE TRAN tdfallA TRIG v(A)  VAL='0.5*VDD' FALL=1 TARG v(Y) VAL='0.5*VDD' FALL=1
.MEASURE TRAN tdriseB TRIG v(B)  VAL='0.5*VDD' RISE=1 TARG v(Y) VAL='0.5*VDD' RISE=1
.MEASURE TRAN tdfallB TRIG v(B)  VAL='0.5*VDD' FALL=1 TARG v(Y) VAL='0.5*VDD' FALL=1
.MEASURE TRAN tdriseC TRIG v(C)  VAL='0.5*VDD' RISE=1 TARG v(Y) VAL='0.5*VDD' RISE=1
.MEASURE TRAN tdfallC TRIG v(C)  VAL='0.5*VDD' FALL=1 TARG v(Y) VAL='0.5*VDD' FALL=1

.MEASURE TRAN Iavg AVG v(Y) FROM=0 TO=10n


.control
save all
op
tran 1n 100n
.endc



.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends
.end
