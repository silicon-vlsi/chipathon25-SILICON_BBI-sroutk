VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp12t3v3__nand3_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__nand3_1 ;
  ORIGIN 0.850 0.000 ;
  SIZE 3.900 BY 8.300 ;
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.850 5.100 3.050 8.300 ;
      LAYER Metal1 ;
        RECT -0.850 7.600 3.050 8.300 ;
        RECT 0.550 6.250 0.800 7.600 ;
        RECT 2.250 5.550 2.500 7.600 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT -0.850 0.000 3.050 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT -0.300 5.450 -0.050 7.250 ;
        RECT 1.400 5.450 1.650 7.250 ;
        RECT -0.300 5.400 1.650 5.450 ;
        RECT -0.300 5.200 1.750 5.400 ;
        RECT 1.250 5.000 1.750 5.200 ;
        RECT -0.100 4.550 0.300 4.950 ;
        RECT 1.400 3.500 1.650 5.000 ;
        RECT 1.900 3.500 2.300 3.950 ;
        RECT -0.300 3.250 1.650 3.500 ;
        RECT -0.300 1.050 -0.050 3.250 ;
        RECT 0.750 2.150 1.150 2.550 ;
      LAYER Metal2 ;
        RECT 1.300 5.000 1.750 5.400 ;
        RECT -0.100 4.550 0.300 4.950 ;
        RECT 1.900 3.500 2.300 3.950 ;
        RECT 0.750 2.150 1.150 2.550 ;
  END
END gf180mcu_osu_sc_gp12t3v3__nand3_1
END LIBRARY

