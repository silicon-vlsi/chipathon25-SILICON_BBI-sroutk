magic
tech gf180mcuD
magscale 1 10
timestamp 1755538115
<< error_p >>
rect 329 780 330 781
rect 359 780 360 781
rect 330 779 331 780
rect 360 779 361 780
<< nwell >>
rect -230 630 980 1270
<< nmos >>
rect -10 210 50 380
rect 160 210 220 380
rect 330 210 390 380
rect 500 210 560 380
rect 680 210 740 380
<< pmos >>
rect 0 720 60 1060
rect 160 720 220 1060
rect 270 780 330 1060
rect 270 720 360 780
rect 500 720 560 1060
rect 690 720 750 1060
<< ndiff >>
rect -110 360 -10 380
rect -110 230 -90 360
rect -40 230 -10 360
rect -110 210 -10 230
rect 50 290 160 380
rect 50 230 80 290
rect 130 230 160 290
rect 50 210 160 230
rect 220 340 330 380
rect 220 230 250 340
rect 300 230 330 340
rect 220 210 330 230
rect 390 290 500 380
rect 390 230 420 290
rect 470 230 500 290
rect 390 210 500 230
rect 560 360 680 380
rect 560 230 590 360
rect 640 230 680 360
rect 560 210 680 230
rect 740 290 840 380
rect 740 230 770 290
rect 820 230 840 290
rect 740 210 840 230
<< pdiff >>
rect -120 1010 0 1060
rect -120 850 -90 1010
rect -40 850 0 1010
rect -120 720 0 850
rect 60 720 160 1060
rect 220 720 270 1060
rect 330 1040 500 1060
rect 330 900 390 1040
rect 470 900 500 1040
rect 330 780 500 900
rect 360 720 500 780
rect 560 1040 690 1060
rect 560 900 590 1040
rect 640 900 690 1040
rect 560 720 690 900
rect 750 1040 870 1060
rect 750 900 780 1040
rect 830 900 870 1040
rect 750 720 870 900
<< ndiffc >>
rect -90 230 -40 360
rect 80 230 130 290
rect 250 230 300 340
rect 420 230 470 290
rect 590 230 640 360
rect 770 230 820 290
<< pdiffc >>
rect -90 850 -40 1010
rect 390 900 470 1040
rect 590 900 640 1040
rect 780 900 830 1040
<< psubdiff >>
rect -180 120 -30 140
rect -180 70 -130 120
rect -80 70 -30 120
rect -180 50 -30 70
rect 60 120 210 140
rect 60 70 110 120
rect 160 70 210 120
rect 60 50 210 70
rect 300 120 450 140
rect 300 70 350 120
rect 400 70 450 120
rect 300 50 450 70
rect 540 120 690 140
rect 540 70 590 120
rect 640 70 690 120
rect 540 50 690 70
rect 780 120 930 140
rect 780 70 820 120
rect 870 70 930 120
rect 780 50 930 70
<< nsubdiff >>
rect -180 1200 -30 1220
rect -180 1150 -130 1200
rect -80 1150 -30 1200
rect -180 1130 -30 1150
rect 60 1200 210 1220
rect 60 1150 110 1200
rect 160 1150 210 1200
rect 60 1130 210 1150
rect 300 1200 450 1220
rect 300 1150 350 1200
rect 400 1150 450 1200
rect 300 1130 450 1150
rect 540 1200 690 1220
rect 540 1150 590 1200
rect 640 1150 690 1200
rect 540 1130 690 1150
rect 780 1200 930 1220
rect 780 1150 830 1200
rect 880 1150 930 1200
rect 780 1130 930 1150
<< psubdiffcont >>
rect -130 70 -80 120
rect 110 70 160 120
rect 350 70 400 120
rect 590 70 640 120
rect 820 70 870 120
<< nsubdiffcont >>
rect -130 1150 -80 1200
rect 110 1150 160 1200
rect 350 1150 400 1200
rect 590 1150 640 1200
rect 830 1150 880 1200
<< polysilicon >>
rect 0 1060 60 1110
rect 160 1060 220 1110
rect 270 1060 330 1110
rect 500 1060 560 1110
rect 690 1060 750 1110
rect 0 670 60 720
rect 10 650 110 670
rect 10 590 30 650
rect 90 590 110 650
rect 10 580 110 590
rect -10 570 110 580
rect -10 380 50 570
rect 160 540 220 720
rect 270 700 360 720
rect 270 670 390 700
rect 500 690 560 720
rect 690 690 750 720
rect 270 650 430 670
rect 330 590 350 650
rect 410 590 430 650
rect 330 570 430 590
rect 500 630 750 690
rect 160 520 280 540
rect 160 460 200 520
rect 260 460 280 520
rect 160 440 280 460
rect 160 380 220 440
rect 330 380 390 570
rect 500 540 560 630
rect 500 520 600 540
rect 500 460 520 520
rect 580 460 600 520
rect 690 460 740 630
rect 500 400 740 460
rect 500 380 560 400
rect 680 380 740 400
rect -10 160 50 210
rect 160 160 220 210
rect 330 160 390 210
rect 500 160 560 210
rect 680 160 740 210
<< polycontact >>
rect 30 590 90 650
rect 350 590 410 650
rect 200 460 260 520
rect 520 460 580 520
<< metal1 >>
rect -210 1200 960 1270
rect -210 1150 -130 1200
rect -80 1150 110 1200
rect 160 1150 350 1200
rect 400 1150 590 1200
rect 640 1150 830 1200
rect 880 1150 960 1200
rect -210 1130 960 1150
rect -90 1010 -40 1060
rect 390 1040 470 1130
rect 390 880 470 900
rect 590 1040 640 1060
rect -90 410 -40 850
rect 590 780 640 900
rect 780 1040 830 1130
rect 780 880 830 900
rect 590 720 610 780
rect 670 720 690 780
rect 10 590 30 650
rect 90 590 110 650
rect 330 590 350 650
rect 410 590 430 650
rect 180 460 200 520
rect 260 460 280 520
rect 490 460 520 520
rect 580 460 600 520
rect 490 420 560 460
rect 490 410 540 420
rect -90 360 540 410
rect 590 370 640 380
rect 590 360 610 370
rect 250 340 300 360
rect -90 210 -40 230
rect 80 290 130 310
rect 80 140 130 230
rect 670 310 690 370
rect 250 210 300 230
rect 420 290 470 310
rect 420 140 470 230
rect 590 210 640 230
rect 770 290 820 310
rect 770 140 820 230
rect -210 120 960 140
rect -210 70 -130 120
rect -80 70 110 120
rect 160 70 350 120
rect 400 70 590 120
rect 640 70 820 120
rect 870 70 960 120
rect -210 0 960 70
<< via1 >>
rect 610 720 670 780
rect 30 590 90 650
rect 350 590 410 650
rect 200 460 260 520
rect 610 360 670 370
rect 610 310 640 360
rect 640 310 670 360
<< metal2 >>
rect 590 780 690 790
rect 590 720 610 780
rect 670 720 690 780
rect 590 710 690 720
rect 10 650 110 660
rect 10 590 30 650
rect 90 590 110 650
rect 10 580 110 590
rect 330 650 430 660
rect 330 590 350 650
rect 410 590 430 650
rect 330 580 430 590
rect 180 520 280 530
rect 180 460 200 520
rect 260 460 280 520
rect 180 450 280 460
rect 610 380 670 710
rect 590 370 690 380
rect 590 310 610 370
rect 670 310 690 370
rect 590 300 690 310
<< labels >>
rlabel metal2 230 490 230 490 1 A
port 1 n
rlabel metal2 380 620 380 620 1 B
port 2 n
rlabel psubdiffcont 130 90 130 90 1 VSS
port 5 n
rlabel via1 640 750 640 750 1 Y
port 3 n
rlabel nsubdiffcont 130 1170 130 1170 1 VDD
port 4 n
flabel metal1 90 1250 540 1260 5 FreeSans 480 0 0 0 VDD
flabel metal1 100 10 550 20 1 FreeSans 480 0 0 0 VSS
flabel polysilicon 200 520 270 540 5 FreeSans 480 0 0 0 B
flabel metal2 620 560 670 590 5 FreeSans 480 0 0 0 Y
flabel polysilicon 40 660 80 670 5 FreeSans 480 0 0 0 C
flabel polysilicon 360 650 420 670 5 FreeSans 480 0 0 0 A
<< end >>
