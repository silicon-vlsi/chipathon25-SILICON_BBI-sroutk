** sch_path: /foss/designs/work/9t_and3_1/gf180mcu_osu_sc_gp9t3v3__and3_1.sch
.subckt gf180mcu_osu_sc_gp9t3v3__and3_1 A B Y C VDD VSS
*.PININFO A:I B:I Y:O C:I VDD:B VSS:B
X1 net1 A VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X0 net1 B VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X2 net1 A net2 VSS nfet_03v3 w=0.85u l=0.3u m=1
X3 net2 B net3 VSS nfet_03v3 w=0.85u l=0.3u m=1
X4 Y net1 VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X5 Y net1 VSS VSS nfet_03v3 w=0.85u l=0.3u m=1
X6 net1 C VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X7 net3 C VSS VSS nfet_03v3 w=0.85u l=0.3u m=1
.ends
