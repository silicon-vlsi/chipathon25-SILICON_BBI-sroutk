VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp12t3v3__and3_1
  CLASS CORE ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__and3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 8.300 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 3.600 1.100 3.900 ;
      LAYER Metal2 ;
        RECT 0.600 3.550 1.100 3.950 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.900 2.950 2.400 3.250 ;
      LAYER Metal2 ;
        RECT 1.900 2.900 2.400 3.300 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.250 5.200 3.700 5.250 ;
        RECT 3.950 5.200 4.200 7.250 ;
        RECT 3.250 4.900 4.200 5.200 ;
        RECT 3.250 4.850 3.700 4.900 ;
        RECT 3.950 1.050 4.200 4.900 ;
      LAYER Metal2 ;
        RECT 3.300 4.850 3.700 5.250 ;
    END
  END Y
  PIN C
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.600 2.300 3.100 2.600 ;
      LAYER Metal2 ;
        RECT 2.600 2.250 3.100 2.650 ;
    END
  END C
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.050 4.800 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 4.800 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 3.100 5.550 3.350 7.600 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 0.000 0.000 4.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 4.550 0.800 7.250 ;
        RECT 2.250 4.550 2.500 7.250 ;
        RECT 3.350 4.550 3.700 4.600 ;
        RECT 0.550 4.250 3.700 4.550 ;
        RECT 1.400 2.250 1.650 4.250 ;
        RECT 3.350 4.200 3.700 4.250 ;
        RECT 0.550 2.000 1.650 2.250 ;
        RECT 0.550 1.050 0.800 2.000 ;
  END
END gf180mcu_osu_sc_gp12t3v3__and3_1
END LIBRARY

