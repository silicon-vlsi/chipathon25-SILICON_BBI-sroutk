magic
tech gf180mcuD
timestamp 1755251668
<< nwell >>
rect 0 102 80 166
<< nmos >>
rect 16 21 22 38
rect 33 21 39 38
rect 52 21 58 38
<< pmos >>
rect 19 111 25 145
rect 30 111 36 145
rect 49 111 55 145
<< ndiff >>
rect 6 36 16 38
rect 6 23 8 36
rect 13 23 16 36
rect 6 21 16 23
rect 22 36 33 38
rect 22 23 25 36
rect 30 23 33 36
rect 22 21 33 23
rect 39 36 52 38
rect 39 23 42 36
rect 47 23 52 36
rect 39 21 52 23
rect 58 36 77 38
rect 58 23 70 36
rect 75 23 77 36
rect 58 21 77 23
<< pdiff >>
rect 9 143 19 145
rect 9 113 11 143
rect 16 113 19 143
rect 9 111 19 113
rect 25 111 30 145
rect 36 111 49 145
rect 55 143 71 145
rect 55 113 58 143
rect 63 113 71 143
rect 55 111 71 113
<< ndiffc >>
rect 8 23 13 36
rect 25 23 30 36
rect 42 23 47 36
rect 70 23 75 36
<< pdiffc >>
rect 11 113 16 143
rect 58 113 63 143
<< psubdiff >>
rect 6 12 21 14
rect 6 7 11 12
rect 16 7 21 12
rect 6 5 21 7
rect 30 12 45 14
rect 30 7 35 12
rect 40 7 45 12
rect 30 5 45 7
rect 54 12 69 14
rect 54 7 59 12
rect 64 7 69 12
rect 54 5 69 7
<< nsubdiff >>
rect 6 159 21 161
rect 6 154 11 159
rect 16 154 21 159
rect 6 152 21 154
rect 30 159 45 161
rect 30 154 35 159
rect 40 154 45 159
rect 30 152 45 154
rect 54 159 69 161
rect 54 154 59 159
rect 64 154 69 159
rect 54 152 69 154
<< psubdiffcont >>
rect 11 7 16 12
rect 35 7 40 12
rect 59 7 64 12
<< nsubdiffcont >>
rect 11 154 16 159
rect 35 154 40 159
rect 59 154 64 159
<< polysilicon >>
rect 19 145 25 150
rect 30 145 36 150
rect 49 145 55 150
rect 19 107 25 111
rect 16 102 25 107
rect 30 108 36 111
rect 49 108 55 111
rect 30 102 39 108
rect 49 102 58 108
rect 16 80 22 102
rect 8 78 22 80
rect 8 72 11 78
rect 17 72 22 78
rect 8 70 22 72
rect 16 38 22 70
rect 33 67 39 102
rect 52 92 58 102
rect 52 90 66 92
rect 52 84 57 90
rect 63 84 66 90
rect 52 82 66 84
rect 33 65 47 67
rect 33 59 39 65
rect 45 59 47 65
rect 33 57 47 59
rect 33 38 39 57
rect 52 38 58 82
rect 16 16 22 21
rect 33 16 39 21
rect 52 16 58 21
<< polycontact >>
rect 11 72 17 78
rect 57 84 63 90
rect 39 59 45 65
<< metal1 >>
rect 0 159 80 166
rect 0 154 11 159
rect 16 154 35 159
rect 40 154 59 159
rect 64 154 80 159
rect 0 152 80 154
rect 11 143 16 152
rect 11 111 16 113
rect 58 143 63 145
rect 58 101 63 113
rect 58 96 75 101
rect 55 84 57 90
rect 63 84 65 90
rect 9 72 11 78
rect 17 72 19 78
rect 70 66 75 96
rect 37 59 39 65
rect 45 59 47 65
rect 68 60 70 66
rect 76 60 78 66
rect 70 50 75 60
rect 25 45 75 50
rect 8 36 13 38
rect 8 14 13 23
rect 25 36 30 45
rect 25 21 30 23
rect 42 36 47 38
rect 42 14 47 23
rect 70 36 75 45
rect 70 21 75 23
rect 0 12 83 14
rect 0 7 11 12
rect 16 7 35 12
rect 40 7 59 12
rect 64 7 83 12
rect 0 0 83 7
<< via1 >>
rect 57 84 63 90
rect 11 72 17 78
rect 39 59 45 65
rect 70 60 76 66
<< metal2 >>
rect 55 90 65 91
rect 55 84 57 90
rect 63 84 65 90
rect 55 83 65 84
rect 9 78 19 79
rect 9 72 11 78
rect 17 72 19 78
rect 9 71 19 72
rect 68 66 78 67
rect 37 65 47 66
rect 37 59 39 65
rect 45 59 47 65
rect 68 60 70 66
rect 76 60 78 66
rect 68 59 78 60
rect 37 58 47 59
<< labels >>
rlabel metal2 14 75 14 75 1 A
port 1 n
rlabel metal2 42 62 42 62 1 B
port 2 n
rlabel nsubdiffcont 14 157 14 157 1 VDD
port 4 n
rlabel psubdiffcont 13 9 13 9 1 VSS
port 5 n
<< end >>
