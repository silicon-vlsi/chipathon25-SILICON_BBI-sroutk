** sch_path: /foss/designs/work/xschem/TB_nand1_3.sch
**.subckt TB_nand1_3

.PARAM PAR_VDD=3.3
.PARAM PAR_CLOAD=5f
.PARAM PAR_SLEW=100p
.PARAM PAR_PER=10n
.CSPARAM PAR_TSTOP='4*PAR_PER'

.INCLUDE ../../core_digital/gf180mcu_osu_sc_gp12t3v3/cells/nand3/gf180mcu_osu_sc_gp12t3v3__nand3_1.spice

**netlist
Xnand 	A B Y C VDD VSS gf180mcu_osu_sc_gp12t3v3__nand3_1
Cload   Y     	VSS  	'PAR_CLOAD' 

**Sources
Vdc   	VDD   	VSS   	PAR_VDD	
VinA   	A    	VSS   	0 	PULSE(0 PAR_VDD '0.1*PAR_PER' PAR_SLEW PAR_SLEW '0.5*PAR_PER' '1.0*PAR_PER')
VinB   	B    	VSS   	0	PULSE(0 PAR_VDD '0.1*PAR_PER' PAR_SLEW PAR_SLEW '1.0*PAR_PER' '2.0*PAR_PER')
VinC   	C    	VSS   	0	PULSE(0 PAR_VDD '0.1*PAR_PER' PAR_SLEW PAR_SLEW '2.0*PAR_PER' '4.0*PAR_PER')
Vgnd	VSS	0	0	

** Rise/Fall 10-90%
.MEASURE TRAN tr1090 TRIG v(Y) VAL='0.1*PAR_VDD' RISE=1 TARG v(Y) VAL='0.9*PAR_VDD' RISE=1
.MEASURE TRAN tf9010 TRIG v(Y) VAL='0.9*PAR_VDD' FALL=1 TARG v(Y) VAL='0.1*PAR_VDD' FALL=1

** Delay Rise Fall
.MEASURE TRAN tdrise TRIG v(A)  VAL='0.5*PAR_VDD' FALL=1 TARG v(Y) VAL='0.5*PAR_VDD' RISE=1
.MEASURE TRAN tdfall TRIG v(A)  VAL='0.5*PAR_VDD' RISE=1 TARG v(Y) VAL='0.5*PAR_VDD' FALL=1

.PLOT v(Y)
.control
save all
op
tran 1p 40n 
.endc



.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends
.end
