* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__and3_2.ext - technology: gf180mcuD

.subckt and3 A B Y C VDD VSS
X0 VDD a_n90_210# Y VDD pfet_03v3 ad=0.561p pd=2.7u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=37400,900
X1 a_250_210# C a_80_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X2 a_n90_210# C VDD VDD pfet_03v3 ad=0.62333p pd=3u as=0.561p ps=2.7u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X3 VSS B a_250_210# VSS nfet_03v3 ad=0.31167p pd=1.86667u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X4 VDD B a_n90_210# VDD pfet_03v3 ad=0.561p pd=2.7u as=0.62333p ps=3u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X5 Y a_n90_210# VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.31167p ps=1.86667u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X6 a_80_210# A a_n90_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.4675p ps=2.8u w=0.85u l=0.3u
**devattr s=18700,560 d=9350,280
X7 Y a_n90_210# VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.561p ps=2.7u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X8 VSS a_n90_210# Y VSS nfet_03v3 ad=0.31167p pd=1.86667u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=18700,560
X9 VDD A a_n90_210# VDD pfet_03v3 ad=0.561p pd=2.7u as=0.62333p ps=3u w=1.7u l=0.3u
**devattr s=37400,900 d=18700,450
.ends

