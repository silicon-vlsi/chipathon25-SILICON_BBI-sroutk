** sch_path: /foss/designs/work/xschem/tb_gf180mcu_osu_sc_gp9t3v3__and3_2.sch
**.subckt tb_gf180mcu_osu_sc_gp9t3v3__and3_2
**** begin user architecture code



** Testbench for AND3_2X

** Parameters
.PARAM VDD=3.3
.PARAM VSS=0
.PARAM CLOAD=50f
.PARAM SLEW=1p

** AND3_2X Design
.INCLUDE gf180mcu_osu_sc_gp9t3v3__and3_2.spice

** Instantiate AND3_2X
Xand A B Y C VDD VDD VDD VDD VSS VSS gf180mcu_osu_sc_gp9t3v3__and3_2

** Load
Cl 	Y	VSS	CLOAD




** Sources
Vdc	VDD	VSS	3.3
Vgnd	VSS	0	0
VinA	A 	VSS	0	PULSE(0 3.3 0 SLEW SLEW 10n 20n)
VinB	B 	VSS	0	PULSE(0 3.3 2n SLEW SLEW 20n 40n)
VinC	C 	VSS	0	PULSE(0 3.3 4n SLEW SLEW 50n 100n)



** Rise/Fall 10-90%
.MEASURE TRAN tr1090 TRIG v(Y) VAL='0.1*VDD' RISE=1 TARG v(Y) VAL='0.9*VDD' RISE=1
.MEASURE TRAN tf9010 TRIG v(Y) VAL='0.9*VDD' FALL=1 TARG v(Y) VAL='0.1*VDD' FALL=1

** Delay Rise Fall
.MEASURE TRAN tdriseA TRIG v(A)  VAL='0.5*VDD' RISE=1 TARG v(Y) VAL='0.5*VDD' RISE=1
.MEASURE TRAN tdfallA TRIG v(A)  VAL='0.5*VDD' RISE=1 TARG v(Y) VAL='0.5*VDD' RISE=1
.MEASURE TRAN tdriseB TRIG v(B)  VAL='0.5*VDD' RISE=1 TARG v(Y) VAL='0.5*VDD' RISE=1
.MEASURE TRAN tdfallB TRIG v(B)  VAL='0.5*VDD' FALL=1 TARG v(Y) VAL='0.5*VDD' FALL=1
.MEASURE TRAN tdriseC TRIG v(C)  VAL='0.5*VDD' RISE=1 TARG v(Y) VAL='0.5*VDD' RISE=1
.MEASURE TRAN tdfallC TRIG v(C)  VAL='0.5*VDD' FALL=1 TARG v(Y) VAL='0.5*VDD' FALL=1

.MEASURE TRAN Iavg AVG Y FROM=0 TO=10n

.control
save all
op
tran 1n 100n
plot v(Y) v(A) v(B) v(C)
.endc
.end



.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends
.end
