magic
tech gf180mcuD
timestamp 1757013610
<< nwell >>
rect 137 102 232 166
<< pwell >>
rect 137 0 232 102
<< nmos >>
rect 156 21 162 38
rect 173 21 179 38
rect 190 21 196 38
rect 207 21 213 38
<< pmos >>
rect 156 111 162 145
rect 173 111 179 145
rect 190 111 196 145
rect 207 111 213 145
<< ndiff >>
rect 146 28 156 38
rect 146 23 148 28
rect 153 23 156 28
rect 146 21 156 23
rect 162 28 173 38
rect 162 23 165 28
rect 170 23 173 28
rect 162 21 173 23
rect 179 28 190 38
rect 179 23 182 28
rect 187 23 190 28
rect 179 21 190 23
rect 196 28 207 38
rect 196 23 199 28
rect 204 23 207 28
rect 196 21 207 23
rect 213 28 223 38
rect 213 23 216 28
rect 221 23 223 28
rect 213 21 223 23
<< pdiff >>
rect 146 143 156 145
rect 146 135 148 143
rect 153 135 156 143
rect 146 111 156 135
rect 162 143 173 145
rect 162 135 165 143
rect 170 135 173 143
rect 162 111 173 135
rect 179 143 190 145
rect 179 135 182 143
rect 187 135 190 143
rect 179 111 190 135
rect 196 143 207 145
rect 196 135 199 143
rect 204 135 207 143
rect 196 111 207 135
rect 213 143 223 145
rect 213 135 216 143
rect 221 135 223 143
rect 213 111 223 135
<< ndiffc >>
rect 148 23 153 28
rect 165 23 170 28
rect 182 23 187 28
rect 199 23 204 28
rect 216 23 221 28
<< pdiffc >>
rect 148 135 153 143
rect 165 135 170 143
rect 182 135 187 143
rect 199 135 204 143
rect 216 135 221 143
<< psubdiff >>
rect 146 12 161 14
rect 146 7 151 12
rect 156 7 161 12
rect 146 5 161 7
rect 177 12 192 14
rect 177 7 182 12
rect 187 7 192 12
rect 177 5 192 7
rect 208 12 223 14
rect 208 7 213 12
rect 218 7 223 12
rect 208 5 223 7
<< nsubdiff >>
rect 146 159 161 161
rect 146 154 151 159
rect 156 154 161 159
rect 146 152 161 154
rect 177 159 192 161
rect 177 154 182 159
rect 187 154 192 159
rect 177 152 192 154
rect 208 159 223 161
rect 208 154 213 159
rect 218 154 223 159
rect 208 152 223 154
<< psubdiffcont >>
rect 151 7 156 12
rect 182 7 187 12
rect 213 7 218 12
<< nsubdiffcont >>
rect 151 154 156 159
rect 182 154 187 159
rect 213 154 218 159
<< polysilicon >>
rect 156 145 162 150
rect 173 145 179 150
rect 190 145 196 150
rect 207 145 213 150
rect 156 82 162 111
rect 150 80 162 82
rect 150 74 152 80
rect 158 74 162 80
rect 150 72 162 74
rect 156 38 162 72
rect 173 95 179 111
rect 173 93 185 95
rect 173 87 177 93
rect 183 87 185 93
rect 173 85 185 87
rect 173 38 179 85
rect 190 69 196 111
rect 207 108 213 111
rect 201 106 213 108
rect 201 100 203 106
rect 209 100 213 106
rect 201 98 213 100
rect 190 67 202 69
rect 190 61 194 67
rect 200 61 202 67
rect 190 59 202 61
rect 190 38 196 59
rect 207 38 213 98
rect 156 16 162 21
rect 173 16 179 21
rect 190 16 196 21
rect 207 16 213 21
<< polycontact >>
rect 152 74 158 80
rect 177 87 183 93
rect 203 100 209 106
rect 194 61 200 67
<< metal1 >>
rect 137 159 232 166
rect 137 154 151 159
rect 156 154 182 159
rect 187 154 213 159
rect 218 154 232 159
rect 137 152 232 154
rect 148 143 153 145
rect 148 126 153 135
rect 165 143 170 145
rect 165 131 170 135
rect 182 143 187 145
rect 182 131 187 135
rect 199 143 204 152
rect 199 133 204 135
rect 216 143 221 145
rect 148 121 209 126
rect 150 74 152 80
rect 158 74 160 80
rect 165 44 170 121
rect 203 106 209 121
rect 203 98 209 100
rect 175 87 177 93
rect 183 87 185 93
rect 216 84 221 135
rect 216 78 218 84
rect 224 78 226 84
rect 192 61 194 67
rect 200 61 202 67
rect 148 39 187 44
rect 148 28 153 39
rect 148 21 153 23
rect 165 28 170 30
rect 165 14 170 23
rect 182 28 187 39
rect 182 21 187 23
rect 199 28 204 30
rect 199 14 204 23
rect 216 28 221 78
rect 216 21 221 23
rect 137 12 232 14
rect 137 7 151 12
rect 156 7 182 12
rect 187 7 213 12
rect 218 7 232 12
rect 137 0 232 7
<< via1 >>
rect 152 74 158 80
rect 203 100 209 106
rect 177 87 183 93
rect 218 78 224 84
rect 194 61 200 67
<< metal2 >>
rect 202 106 210 108
rect 202 100 203 106
rect 209 100 210 106
rect 202 98 210 100
rect 175 93 185 94
rect 175 87 177 93
rect 183 87 185 93
rect 175 86 185 87
rect 216 84 226 85
rect 150 80 160 81
rect 150 74 152 80
rect 158 74 160 80
rect 216 78 218 84
rect 224 78 226 84
rect 216 77 226 78
rect 150 73 160 74
rect 192 67 202 68
rect 192 61 194 67
rect 200 61 202 67
rect 192 60 202 61
<< labels >>
flabel metal1 161 155 177 163 0 FreeSans 48 0 0 0 VDD
port 5 nsew
flabel metal1 161 2 177 10 0 FreeSans 48 0 0 0 VSS
port 6 nsew
flabel metal2 192 60 202 68 0 FreeSans 48 0 0 0 A
port 1 nsew
flabel metal2 175 86 185 94 0 FreeSans 48 0 0 0 B
port 2 nsew
flabel metal2 150 73 160 81 0 FreeSans 48 0 0 0 C
port 3 nsew
flabel metal2 216 77 226 85 0 FreeSans 48 0 0 0 Y
port 4 nsew
<< properties >>
string FIXED_BBOX 137 0 232 166
<< end >>
