VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp12t3v3__and3_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__and3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.750 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 3.600 1.100 3.900 ;
      LAYER Metal2 ;
        RECT 0.600 3.550 1.100 3.950 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.900 2.950 2.400 3.250 ;
      LAYER Metal2 ;
        RECT 1.900 2.900 2.400 3.300 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.950 5.300 4.200 7.250 ;
        RECT 3.950 4.900 4.400 5.300 ;
        RECT 3.950 1.050 4.200 4.900 ;
      LAYER Metal2 ;
        RECT 3.950 4.900 4.400 5.300 ;
    END
  END Y
  PIN C
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.700 2.300 3.200 2.600 ;
      LAYER Metal2 ;
        RECT 2.700 2.250 3.200 2.650 ;
    END
  END C
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 4.750 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 4.750 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 3.100 5.550 3.350 7.600 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.000 0.000 4.750 5.100 ;
      LAYER Metal1 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 0.000 0.000 4.750 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 4.600 0.800 7.250 ;
        RECT 2.250 4.600 2.500 7.250 ;
        RECT 0.550 4.300 3.700 4.600 ;
        RECT 1.400 2.250 1.650 4.300 ;
        RECT 0.550 2.000 1.650 2.250 ;
        RECT 0.550 1.050 0.800 2.000 ;
  END
END gf180mcu_osu_sc_gp12t3v3__and3_1
END LIBRARY

