** sch_path: /foss/designs/work/9tnand3/gf180mcu_osu_sc_gp9t3v3__nand3_1.sch
.subckt gf180mcu_osu_sc_gp9t3v3__nand3_1 A B Y C VDD VSS
*.PININFO A:I B:I Y:O C:I VDD:B VSS:B
X1 Y A VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X0 Y B VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
X2 Y A net1 VSS nfet_03v3 w=0.85u l=0.3u m=1
X3 net1 B net2 VSS nfet_03v3 w=0.85u l=0.3u m=1
X4 net2 C VSS VSS nfet_03v3 w=0.85u l=0.3u m=1
X5 Y C VDD VDD pfet_03v3 w=1.7u l=0.3u m=1
.ends
