** sch_path: /foss/designs/work/9t_nand3/tb_gf180mcu_osu_sc_gp9t3v3__nand3_1.sch
**.subckt tb_gf180mcu_osu_sc_gp9t3v3__nand3_1
**** begin user architecture code


.PARAM PAR_VDD=3.3
.CSPARAM CPAR_VDD=PAR_VDD
.PARAM PAR_CLOAD=50f
.PARAM PAR_SLEW=100p
.PARAM PAR_PER=10n
.CSPARAM CPAR_PER=PAR_PER
.PARAM PAR_DEL='0.1*PAR_PER'
.CSPARAM CPAR_DEL=PAR_DEL

.INCLUDE gf180mcu_osu_sc_gp9t3v3__nand3_1.spice

**netlist
Xor3 A B Y C VDD VSS gf180mcu_osu_sc_gp9t3v3__nand3_1
Cload   Y     	VSS  	'PAR_CLOAD'

**Sources
Vdc   	VDD   	VSS   	PAR_VDD
VinA   	A    	VSS   	0 	PULSE( 'PAR_VDD' 0 PAR_DEL PAR_SLEW PAR_SLEW '0.5*PAR_PER' '1.0*PAR_PER')
VinB   	B    	VSS   	0	PULSE( 'PAR_VDD' 0 PAR_DEL PAR_SLEW PAR_SLEW '1.0*PAR_PER' '2.0*PAR_PER')
VinC   	C    	VSS   	0	PULSE( 'PAR_VDD' 0 PAR_DEL PAR_SLEW PAR_SLEW '2.0*PAR_PER' '4.0*PAR_PER')
Vgnd	VSS	0	0

** Rise/Fall 10-90%
.MEASURE TRAN tr1090 TRIG v(Y) VAL='0.1*PAR_VDD' RISE=1 TARG v(Y) VAL='0.9*PAR_VDD' RISE=1
.MEASURE TRAN tf9010 TRIG v(Y) VAL='0.9*PAR_VDD' FALL=1 TARG v(Y) VAL='0.1*PAR_VDD' FALL=1

** Delay Rise Fall
.MEASURE TRAN tdrise TRIG v(A)  VAL='0.5*PAR_VDD' RISE=1 TARG v(Y) VAL='0.5*PAR_VDD' RISE=1
.MEASURE TRAN tdfall TRIG v(A)  VAL='0.5*PAR_VDD' FALL=1 TARG v(Y) VAL='0.5*PAR_VDD' FALL=1

**Leakage current and average current
.MEASURE TRAN iavg AVG vdc#branch FROM=PAR_DEL TO='PAR_DEL+PAR_PER'
.MEASURE TRAN ileak AVG vdc#branch FROM='PAR_DEL+0.4*PAR_PER' TO='PAR_DEL+0.45*PAR_PER'

.control
save all
OP
TRAN 1p 41n

PLOT v(Y) 'CPAR_VDD + v(A)' '2*CPAR_VDD + v(B)' '3*CPAR_VDD + v(C)'
LET cut-tstart=CPAR_DEL
LET cut-tstop='0.75*CPAR_PER'
cutout
PLOT v(Y) v(A)

.endc




.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends
.end
