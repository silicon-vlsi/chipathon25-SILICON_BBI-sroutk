magic
tech gf180mcuD
magscale 1 10
timestamp 1755791114
<< error_p >>
rect 1250 899 1261 900
rect 1289 899 1300 900
<< nwell >>
rect 1140 630 1920 1270
<< nmos >>
rect 1330 210 1390 380
rect 1500 210 1560 380
rect 1670 210 1730 380
<< pmos >>
rect 1330 720 1390 1060
rect 1500 720 1560 1060
rect 1670 720 1730 1060
<< ndiff >>
rect 1230 280 1330 380
rect 1230 230 1250 280
rect 1300 230 1330 280
rect 1230 210 1330 230
rect 1390 280 1500 380
rect 1390 230 1420 280
rect 1470 230 1500 280
rect 1390 210 1500 230
rect 1560 280 1670 380
rect 1560 230 1590 280
rect 1640 230 1670 280
rect 1560 210 1670 230
rect 1730 280 1830 380
rect 1730 230 1760 280
rect 1810 230 1830 280
rect 1730 210 1830 230
<< pdiff >>
rect 1230 1040 1330 1060
rect 1230 910 1250 1040
rect 1300 910 1330 1040
rect 1230 720 1330 910
rect 1390 1040 1500 1060
rect 1390 910 1420 1040
rect 1470 910 1500 1040
rect 1390 720 1500 910
rect 1560 1040 1670 1060
rect 1560 910 1590 1040
rect 1640 910 1670 1040
rect 1560 720 1670 910
rect 1730 1040 1830 1060
rect 1730 910 1760 1040
rect 1810 910 1830 1040
rect 1730 720 1830 910
<< ndiffc >>
rect 1250 230 1300 280
rect 1420 230 1470 280
rect 1590 230 1640 280
rect 1760 230 1810 280
<< pdiffc >>
rect 1250 910 1300 1040
rect 1420 910 1470 1040
rect 1590 910 1640 1040
rect 1760 910 1810 1040
<< psubdiff >>
rect 1230 120 1380 140
rect 1230 70 1280 120
rect 1330 70 1380 120
rect 1230 50 1380 70
rect 1680 120 1830 140
rect 1680 70 1730 120
rect 1780 70 1830 120
rect 1680 50 1830 70
<< nsubdiff >>
rect 1230 1200 1380 1220
rect 1230 1150 1280 1200
rect 1330 1150 1380 1200
rect 1230 1130 1380 1150
rect 1680 1200 1830 1220
rect 1680 1150 1730 1200
rect 1780 1150 1830 1200
rect 1680 1130 1830 1150
<< psubdiffcont >>
rect 1280 70 1330 120
rect 1730 70 1780 120
<< nsubdiffcont >>
rect 1280 1150 1330 1200
rect 1730 1150 1780 1200
<< polysilicon >>
rect 1330 1060 1390 1110
rect 1500 1060 1560 1110
rect 1670 1060 1730 1110
rect 1330 510 1390 720
rect 1270 490 1390 510
rect 1270 430 1290 490
rect 1350 430 1390 490
rect 1270 410 1390 430
rect 1330 380 1390 410
rect 1500 510 1560 720
rect 1670 700 1730 720
rect 1610 680 1730 700
rect 1610 620 1630 680
rect 1690 620 1730 680
rect 1610 600 1730 620
rect 1500 490 1620 510
rect 1500 430 1540 490
rect 1600 430 1620 490
rect 1500 410 1620 430
rect 1500 380 1560 410
rect 1670 380 1730 600
rect 1330 160 1390 210
rect 1500 160 1560 210
rect 1670 160 1730 210
<< polycontact >>
rect 1290 430 1350 490
rect 1630 620 1690 680
rect 1540 430 1600 490
<< metal1 >>
rect 1140 1200 1920 1270
rect 1140 1150 1280 1200
rect 1330 1150 1730 1200
rect 1780 1150 1920 1200
rect 1140 1130 1920 1150
rect 1250 1040 1300 1130
rect 1250 900 1300 910
rect 1420 1040 1470 1060
rect 1420 890 1470 910
rect 1590 1040 1640 1060
rect 1590 890 1640 910
rect 1760 1040 1810 1060
rect 1760 830 1810 910
rect 1420 780 1810 830
rect 1270 430 1290 490
rect 1350 430 1370 490
rect 1250 280 1300 300
rect 1250 140 1300 230
rect 1420 280 1470 780
rect 1610 620 1630 680
rect 1690 620 1710 680
rect 1760 490 1810 780
rect 1520 430 1540 490
rect 1600 430 1620 490
rect 1760 430 1830 490
rect 1890 430 1910 490
rect 1420 210 1470 230
rect 1590 280 1640 300
rect 1590 140 1640 230
rect 1760 280 1810 430
rect 1760 210 1810 230
rect 1140 120 1920 140
rect 1140 70 1280 120
rect 1330 70 1730 120
rect 1780 70 1920 120
rect 1140 0 1920 70
<< via1 >>
rect 1290 430 1350 490
rect 1630 620 1690 680
rect 1540 430 1600 490
rect 1830 430 1890 490
<< metal2 >>
rect 1610 680 1710 690
rect 1610 620 1630 680
rect 1690 620 1710 680
rect 1610 610 1710 620
rect 1270 490 1370 500
rect 1270 430 1290 490
rect 1350 430 1370 490
rect 1270 420 1370 430
rect 1520 490 1620 500
rect 1520 430 1540 490
rect 1600 430 1620 490
rect 1520 420 1620 430
rect 1810 490 1910 500
rect 1810 430 1830 490
rect 1890 430 1910 490
rect 1810 420 1910 430
<< labels >>
flabel metal2 1290 430 1350 490 0 FreeSans 480 0 0 0 A
flabel metal2 1540 430 1600 490 0 FreeSans 480 0 0 0 B
flabel metal2 1630 620 1690 680 0 FreeSans 480 0 0 0 C
flabel via1 1830 430 1890 490 0 FreeSans 480 0 0 0 Y
flabel metal1 1150 1210 1240 1250 0 FreeSans 320 0 0 0 VDD
flabel metal1 1140 20 1230 60 0 FreeSans 320 0 0 0 VSS
rlabel pdiffc 1250 910 1300 1040 1 net1
rlabel ndiffc 1250 230 1300 280 1 net2
rlabel ndiffc 1420 230 1470 280 1 net3
<< end >>
