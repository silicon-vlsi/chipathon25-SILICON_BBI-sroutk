* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__and3_2.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__and3_2 A B Y C VDD VSS
X0 VDD a_n90_210# Y VDD pfet_03v3 ad=0.561p pd=2.7u as=0.4675p ps=2.25u w=1.7u l=0.3u
**devattr s=18700,450 d=37400,900
X1 a_250_210# B a_80_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X2 a_n90_210# B VDD VDD pfet_03v3 ad=0.62333p pd=3u as=0.561p ps=2.7u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X3 VSS C a_250_210# VSS nfet_03v3 ad=0.31167p pd=1.86667u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X4 VDD C a_n90_210# VDD pfet_03v3 ad=0.561p pd=2.7u as=0.62333p ps=3u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X5 Y a_n90_210# VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.31167p ps=1.86667u w=0.85u l=0.3u
**devattr s=9350,280 d=9350,280
X6 a_80_210# A a_n90_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.4675p ps=2.8u w=0.85u l=0.3u
**devattr s=18700,560 d=9350,280
X7 Y a_n90_210# VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.561p ps=2.7u w=1.7u l=0.3u
**devattr s=18700,450 d=18700,450
X8 VSS a_n90_210# Y VSS nfet_03v3 ad=0.31167p pd=1.86667u as=0.23375p ps=1.4u w=0.85u l=0.3u
**devattr s=9350,280 d=18700,560
X9 VDD A a_n90_210# VDD pfet_03v3 ad=0.561p pd=2.7u as=0.62333p ps=3u w=1.7u l=0.3u
**devattr s=37400,900 d=18700,450
C0 C Y 0.03198f
C1 VDD A 0.12462f
C2 B a_n90_210# 0.1824f
C3 C a_250_210# 0.02615f
C4 a_n90_210# Y 0.28319f
C5 B A 0.06819f
C6 A a_n90_210# 0.22916f
C7 VDD C 0.08642f
C8 a_n90_210# a_80_210# 0.08029f
C9 B VDD 0.11714f
C10 B C 0.09692f
C11 VDD a_n90_210# 0.6672f
C12 C a_n90_210# 0.14156f
C13 a_80_210# a_250_210# 0.05362f
C14 VDD Y 0.18192f
C15 Y VSS 0.31276f
C16 C VSS 0.32317f
C17 B VSS 0.28589f
C18 A VSS 0.34197f
C19 VDD VSS 2.49623f
C20 a_250_210# VSS 0.08046f
C21 a_80_210# VSS 0.04401f
C22 a_n90_210# VSS 0.83934f
.ends

